module division_LUT_ap_fixed_16_10_s15 #(
)(
    input logic [16-1:0] number_in,
    output logic [16-1:0] reciprocal

);

    logic [32767:0] reciprocal_LUT [16-1:0];

    always_comb begin
        case (number_in[16-1:16-15])
        15'b000000000000001 : reciprocal = 16'b0000001000000000;
        15'b000000000000010 : reciprocal = 16'b0000000100000000;
        15'b000000000000011 : reciprocal = 16'b0000000010101011;
        15'b000000000000100 : reciprocal = 16'b0000000010000000;
        15'b000000000000101 : reciprocal = 16'b0000000001100110;
        15'b000000000000110 : reciprocal = 16'b0000000001010101;
        15'b000000000000111 : reciprocal = 16'b0000000001001001;
        15'b000000000001000 : reciprocal = 16'b0000000001000000;
        15'b000000000001001 : reciprocal = 16'b0000000000111001;
        15'b000000000001010 : reciprocal = 16'b0000000000110011;
        15'b000000000001011 : reciprocal = 16'b0000000000101111;
        15'b000000000001100 : reciprocal = 16'b0000000000101011;
        15'b000000000001101 : reciprocal = 16'b0000000000100111;
        15'b000000000001110 : reciprocal = 16'b0000000000100101;
        15'b000000000001111 : reciprocal = 16'b0000000000100010;
        15'b000000000010000 : reciprocal = 16'b0000000000100000;
        15'b000000000010001 : reciprocal = 16'b0000000000011110;
        15'b000000000010010 : reciprocal = 16'b0000000000011100;
        15'b000000000010011 : reciprocal = 16'b0000000000011011;
        15'b000000000010100 : reciprocal = 16'b0000000000011010;
        15'b000000000010101 : reciprocal = 16'b0000000000011000;
        15'b000000000010110 : reciprocal = 16'b0000000000010111;
        15'b000000000010111 : reciprocal = 16'b0000000000010110;
        15'b000000000011000 : reciprocal = 16'b0000000000010101;
        15'b000000000011001 : reciprocal = 16'b0000000000010100;
        15'b000000000011010 : reciprocal = 16'b0000000000010100;
        15'b000000000011011 : reciprocal = 16'b0000000000010011;
        15'b000000000011100 : reciprocal = 16'b0000000000010010;
        15'b000000000011101 : reciprocal = 16'b0000000000010010;
        15'b000000000011110 : reciprocal = 16'b0000000000010001;
        15'b000000000011111 : reciprocal = 16'b0000000000010001;
        15'b000000000100000 : reciprocal = 16'b0000000000010000;
        15'b000000000100001 : reciprocal = 16'b0000000000010000;
        15'b000000000100010 : reciprocal = 16'b0000000000001111;
        15'b000000000100011 : reciprocal = 16'b0000000000001111;
        15'b000000000100100 : reciprocal = 16'b0000000000001110;
        15'b000000000100101 : reciprocal = 16'b0000000000001110;
        15'b000000000100110 : reciprocal = 16'b0000000000001101;
        15'b000000000100111 : reciprocal = 16'b0000000000001101;
        15'b000000000101000 : reciprocal = 16'b0000000000001101;
        15'b000000000101001 : reciprocal = 16'b0000000000001100;
        15'b000000000101010 : reciprocal = 16'b0000000000001100;
        15'b000000000101011 : reciprocal = 16'b0000000000001100;
        15'b000000000101100 : reciprocal = 16'b0000000000001100;
        15'b000000000101101 : reciprocal = 16'b0000000000001011;
        15'b000000000101110 : reciprocal = 16'b0000000000001011;
        15'b000000000101111 : reciprocal = 16'b0000000000001011;
        15'b000000000110000 : reciprocal = 16'b0000000000001011;
        15'b000000000110001 : reciprocal = 16'b0000000000001010;
        15'b000000000110010 : reciprocal = 16'b0000000000001010;
        15'b000000000110011 : reciprocal = 16'b0000000000001010;
        15'b000000000110100 : reciprocal = 16'b0000000000001010;
        15'b000000000110101 : reciprocal = 16'b0000000000001010;
        15'b000000000110110 : reciprocal = 16'b0000000000001001;
        15'b000000000110111 : reciprocal = 16'b0000000000001001;
        15'b000000000111000 : reciprocal = 16'b0000000000001001;
        15'b000000000111001 : reciprocal = 16'b0000000000001001;
        15'b000000000111010 : reciprocal = 16'b0000000000001001;
        15'b000000000111011 : reciprocal = 16'b0000000000001001;
        15'b000000000111100 : reciprocal = 16'b0000000000001001;
        15'b000000000111101 : reciprocal = 16'b0000000000001000;
        15'b000000000111110 : reciprocal = 16'b0000000000001000;
        15'b000000000111111 : reciprocal = 16'b0000000000001000;
        15'b000000001000000 : reciprocal = 16'b0000000000001000;
        15'b000000001000001 : reciprocal = 16'b0000000000001000;
        15'b000000001000010 : reciprocal = 16'b0000000000001000;
        15'b000000001000011 : reciprocal = 16'b0000000000001000;
        15'b000000001000100 : reciprocal = 16'b0000000000001000;
        15'b000000001000101 : reciprocal = 16'b0000000000000111;
        15'b000000001000110 : reciprocal = 16'b0000000000000111;
        15'b000000001000111 : reciprocal = 16'b0000000000000111;
        15'b000000001001000 : reciprocal = 16'b0000000000000111;
        15'b000000001001001 : reciprocal = 16'b0000000000000111;
        15'b000000001001010 : reciprocal = 16'b0000000000000111;
        15'b000000001001011 : reciprocal = 16'b0000000000000111;
        15'b000000001001100 : reciprocal = 16'b0000000000000111;
        15'b000000001001101 : reciprocal = 16'b0000000000000111;
        15'b000000001001110 : reciprocal = 16'b0000000000000111;
        15'b000000001001111 : reciprocal = 16'b0000000000000110;
        15'b000000001010000 : reciprocal = 16'b0000000000000110;
        15'b000000001010001 : reciprocal = 16'b0000000000000110;
        15'b000000001010010 : reciprocal = 16'b0000000000000110;
        15'b000000001010011 : reciprocal = 16'b0000000000000110;
        15'b000000001010100 : reciprocal = 16'b0000000000000110;
        15'b000000001010101 : reciprocal = 16'b0000000000000110;
        15'b000000001010110 : reciprocal = 16'b0000000000000110;
        15'b000000001010111 : reciprocal = 16'b0000000000000110;
        15'b000000001011000 : reciprocal = 16'b0000000000000110;
        15'b000000001011001 : reciprocal = 16'b0000000000000110;
        15'b000000001011010 : reciprocal = 16'b0000000000000110;
        15'b000000001011011 : reciprocal = 16'b0000000000000110;
        15'b000000001011100 : reciprocal = 16'b0000000000000110;
        15'b000000001011101 : reciprocal = 16'b0000000000000110;
        15'b000000001011110 : reciprocal = 16'b0000000000000101;
        15'b000000001011111 : reciprocal = 16'b0000000000000101;
        15'b000000001100000 : reciprocal = 16'b0000000000000101;
        15'b000000001100001 : reciprocal = 16'b0000000000000101;
        15'b000000001100010 : reciprocal = 16'b0000000000000101;
        15'b000000001100011 : reciprocal = 16'b0000000000000101;
        15'b000000001100100 : reciprocal = 16'b0000000000000101;
        15'b000000001100101 : reciprocal = 16'b0000000000000101;
        15'b000000001100110 : reciprocal = 16'b0000000000000101;
        15'b000000001100111 : reciprocal = 16'b0000000000000101;
        15'b000000001101000 : reciprocal = 16'b0000000000000101;
        15'b000000001101001 : reciprocal = 16'b0000000000000101;
        15'b000000001101010 : reciprocal = 16'b0000000000000101;
        15'b000000001101011 : reciprocal = 16'b0000000000000101;
        15'b000000001101100 : reciprocal = 16'b0000000000000101;
        15'b000000001101101 : reciprocal = 16'b0000000000000101;
        15'b000000001101110 : reciprocal = 16'b0000000000000101;
        15'b000000001101111 : reciprocal = 16'b0000000000000101;
        15'b000000001110000 : reciprocal = 16'b0000000000000101;
        15'b000000001110001 : reciprocal = 16'b0000000000000101;
        15'b000000001110010 : reciprocal = 16'b0000000000000100;
        15'b000000001110011 : reciprocal = 16'b0000000000000100;
        15'b000000001110100 : reciprocal = 16'b0000000000000100;
        15'b000000001110101 : reciprocal = 16'b0000000000000100;
        15'b000000001110110 : reciprocal = 16'b0000000000000100;
        15'b000000001110111 : reciprocal = 16'b0000000000000100;
        15'b000000001111000 : reciprocal = 16'b0000000000000100;
        15'b000000001111001 : reciprocal = 16'b0000000000000100;
        15'b000000001111010 : reciprocal = 16'b0000000000000100;
        15'b000000001111011 : reciprocal = 16'b0000000000000100;
        15'b000000001111100 : reciprocal = 16'b0000000000000100;
        15'b000000001111101 : reciprocal = 16'b0000000000000100;
        15'b000000001111110 : reciprocal = 16'b0000000000000100;
        15'b000000001111111 : reciprocal = 16'b0000000000000100;
        15'b000000010000000 : reciprocal = 16'b0000000000000100;
        15'b000000010000001 : reciprocal = 16'b0000000000000100;
        15'b000000010000010 : reciprocal = 16'b0000000000000100;
        15'b000000010000011 : reciprocal = 16'b0000000000000100;
        15'b000000010000100 : reciprocal = 16'b0000000000000100;
        15'b000000010000101 : reciprocal = 16'b0000000000000100;
        15'b000000010000110 : reciprocal = 16'b0000000000000100;
        15'b000000010000111 : reciprocal = 16'b0000000000000100;
        15'b000000010001000 : reciprocal = 16'b0000000000000100;
        15'b000000010001001 : reciprocal = 16'b0000000000000100;
        15'b000000010001010 : reciprocal = 16'b0000000000000100;
        15'b000000010001011 : reciprocal = 16'b0000000000000100;
        15'b000000010001100 : reciprocal = 16'b0000000000000100;
        15'b000000010001101 : reciprocal = 16'b0000000000000100;
        15'b000000010001110 : reciprocal = 16'b0000000000000100;
        15'b000000010001111 : reciprocal = 16'b0000000000000100;
        15'b000000010010000 : reciprocal = 16'b0000000000000100;
        15'b000000010010001 : reciprocal = 16'b0000000000000100;
        15'b000000010010010 : reciprocal = 16'b0000000000000100;
        15'b000000010010011 : reciprocal = 16'b0000000000000011;
        15'b000000010010100 : reciprocal = 16'b0000000000000011;
        15'b000000010010101 : reciprocal = 16'b0000000000000011;
        15'b000000010010110 : reciprocal = 16'b0000000000000011;
        15'b000000010010111 : reciprocal = 16'b0000000000000011;
        15'b000000010011000 : reciprocal = 16'b0000000000000011;
        15'b000000010011001 : reciprocal = 16'b0000000000000011;
        15'b000000010011010 : reciprocal = 16'b0000000000000011;
        15'b000000010011011 : reciprocal = 16'b0000000000000011;
        15'b000000010011100 : reciprocal = 16'b0000000000000011;
        15'b000000010011101 : reciprocal = 16'b0000000000000011;
        15'b000000010011110 : reciprocal = 16'b0000000000000011;
        15'b000000010011111 : reciprocal = 16'b0000000000000011;
        15'b000000010100000 : reciprocal = 16'b0000000000000011;
        15'b000000010100001 : reciprocal = 16'b0000000000000011;
        15'b000000010100010 : reciprocal = 16'b0000000000000011;
        15'b000000010100011 : reciprocal = 16'b0000000000000011;
        15'b000000010100100 : reciprocal = 16'b0000000000000011;
        15'b000000010100101 : reciprocal = 16'b0000000000000011;
        15'b000000010100110 : reciprocal = 16'b0000000000000011;
        15'b000000010100111 : reciprocal = 16'b0000000000000011;
        15'b000000010101000 : reciprocal = 16'b0000000000000011;
        15'b000000010101001 : reciprocal = 16'b0000000000000011;
        15'b000000010101010 : reciprocal = 16'b0000000000000011;
        15'b000000010101011 : reciprocal = 16'b0000000000000011;
        15'b000000010101100 : reciprocal = 16'b0000000000000011;
        15'b000000010101101 : reciprocal = 16'b0000000000000011;
        15'b000000010101110 : reciprocal = 16'b0000000000000011;
        15'b000000010101111 : reciprocal = 16'b0000000000000011;
        15'b000000010110000 : reciprocal = 16'b0000000000000011;
        15'b000000010110001 : reciprocal = 16'b0000000000000011;
        15'b000000010110010 : reciprocal = 16'b0000000000000011;
        15'b000000010110011 : reciprocal = 16'b0000000000000011;
        15'b000000010110100 : reciprocal = 16'b0000000000000011;
        15'b000000010110101 : reciprocal = 16'b0000000000000011;
        15'b000000010110110 : reciprocal = 16'b0000000000000011;
        15'b000000010110111 : reciprocal = 16'b0000000000000011;
        15'b000000010111000 : reciprocal = 16'b0000000000000011;
        15'b000000010111001 : reciprocal = 16'b0000000000000011;
        15'b000000010111010 : reciprocal = 16'b0000000000000011;
        15'b000000010111011 : reciprocal = 16'b0000000000000011;
        15'b000000010111100 : reciprocal = 16'b0000000000000011;
        15'b000000010111101 : reciprocal = 16'b0000000000000011;
        15'b000000010111110 : reciprocal = 16'b0000000000000011;
        15'b000000010111111 : reciprocal = 16'b0000000000000011;
        15'b000000011000000 : reciprocal = 16'b0000000000000011;
        15'b000000011000001 : reciprocal = 16'b0000000000000011;
        15'b000000011000010 : reciprocal = 16'b0000000000000011;
        15'b000000011000011 : reciprocal = 16'b0000000000000011;
        15'b000000011000100 : reciprocal = 16'b0000000000000011;
        15'b000000011000101 : reciprocal = 16'b0000000000000011;
        15'b000000011000110 : reciprocal = 16'b0000000000000011;
        15'b000000011000111 : reciprocal = 16'b0000000000000011;
        15'b000000011001000 : reciprocal = 16'b0000000000000011;
        15'b000000011001001 : reciprocal = 16'b0000000000000011;
        15'b000000011001010 : reciprocal = 16'b0000000000000011;
        15'b000000011001011 : reciprocal = 16'b0000000000000011;
        15'b000000011001100 : reciprocal = 16'b0000000000000011;
        15'b000000011001101 : reciprocal = 16'b0000000000000010;
        15'b000000011001110 : reciprocal = 16'b0000000000000010;
        15'b000000011001111 : reciprocal = 16'b0000000000000010;
        15'b000000011010000 : reciprocal = 16'b0000000000000010;
        15'b000000011010001 : reciprocal = 16'b0000000000000010;
        15'b000000011010010 : reciprocal = 16'b0000000000000010;
        15'b000000011010011 : reciprocal = 16'b0000000000000010;
        15'b000000011010100 : reciprocal = 16'b0000000000000010;
        15'b000000011010101 : reciprocal = 16'b0000000000000010;
        15'b000000011010110 : reciprocal = 16'b0000000000000010;
        15'b000000011010111 : reciprocal = 16'b0000000000000010;
        15'b000000011011000 : reciprocal = 16'b0000000000000010;
        15'b000000011011001 : reciprocal = 16'b0000000000000010;
        15'b000000011011010 : reciprocal = 16'b0000000000000010;
        15'b000000011011011 : reciprocal = 16'b0000000000000010;
        15'b000000011011100 : reciprocal = 16'b0000000000000010;
        15'b000000011011101 : reciprocal = 16'b0000000000000010;
        15'b000000011011110 : reciprocal = 16'b0000000000000010;
        15'b000000011011111 : reciprocal = 16'b0000000000000010;
        15'b000000011100000 : reciprocal = 16'b0000000000000010;
        15'b000000011100001 : reciprocal = 16'b0000000000000010;
        15'b000000011100010 : reciprocal = 16'b0000000000000010;
        15'b000000011100011 : reciprocal = 16'b0000000000000010;
        15'b000000011100100 : reciprocal = 16'b0000000000000010;
        15'b000000011100101 : reciprocal = 16'b0000000000000010;
        15'b000000011100110 : reciprocal = 16'b0000000000000010;
        15'b000000011100111 : reciprocal = 16'b0000000000000010;
        15'b000000011101000 : reciprocal = 16'b0000000000000010;
        15'b000000011101001 : reciprocal = 16'b0000000000000010;
        15'b000000011101010 : reciprocal = 16'b0000000000000010;
        15'b000000011101011 : reciprocal = 16'b0000000000000010;
        15'b000000011101100 : reciprocal = 16'b0000000000000010;
        15'b000000011101101 : reciprocal = 16'b0000000000000010;
        15'b000000011101110 : reciprocal = 16'b0000000000000010;
        15'b000000011101111 : reciprocal = 16'b0000000000000010;
        15'b000000011110000 : reciprocal = 16'b0000000000000010;
        15'b000000011110001 : reciprocal = 16'b0000000000000010;
        15'b000000011110010 : reciprocal = 16'b0000000000000010;
        15'b000000011110011 : reciprocal = 16'b0000000000000010;
        15'b000000011110100 : reciprocal = 16'b0000000000000010;
        15'b000000011110101 : reciprocal = 16'b0000000000000010;
        15'b000000011110110 : reciprocal = 16'b0000000000000010;
        15'b000000011110111 : reciprocal = 16'b0000000000000010;
        15'b000000011111000 : reciprocal = 16'b0000000000000010;
        15'b000000011111001 : reciprocal = 16'b0000000000000010;
        15'b000000011111010 : reciprocal = 16'b0000000000000010;
        15'b000000011111011 : reciprocal = 16'b0000000000000010;
        15'b000000011111100 : reciprocal = 16'b0000000000000010;
        15'b000000011111101 : reciprocal = 16'b0000000000000010;
        15'b000000011111110 : reciprocal = 16'b0000000000000010;
        15'b000000011111111 : reciprocal = 16'b0000000000000010;
        15'b000000100000000 : reciprocal = 16'b0000000000000010;
        15'b000000100000001 : reciprocal = 16'b0000000000000010;
        15'b000000100000010 : reciprocal = 16'b0000000000000010;
        15'b000000100000011 : reciprocal = 16'b0000000000000010;
        15'b000000100000100 : reciprocal = 16'b0000000000000010;
        15'b000000100000101 : reciprocal = 16'b0000000000000010;
        15'b000000100000110 : reciprocal = 16'b0000000000000010;
        15'b000000100000111 : reciprocal = 16'b0000000000000010;
        15'b000000100001000 : reciprocal = 16'b0000000000000010;
        15'b000000100001001 : reciprocal = 16'b0000000000000010;
        15'b000000100001010 : reciprocal = 16'b0000000000000010;
        15'b000000100001011 : reciprocal = 16'b0000000000000010;
        15'b000000100001100 : reciprocal = 16'b0000000000000010;
        15'b000000100001101 : reciprocal = 16'b0000000000000010;
        15'b000000100001110 : reciprocal = 16'b0000000000000010;
        15'b000000100001111 : reciprocal = 16'b0000000000000010;
        15'b000000100010000 : reciprocal = 16'b0000000000000010;
        15'b000000100010001 : reciprocal = 16'b0000000000000010;
        15'b000000100010010 : reciprocal = 16'b0000000000000010;
        15'b000000100010011 : reciprocal = 16'b0000000000000010;
        15'b000000100010100 : reciprocal = 16'b0000000000000010;
        15'b000000100010101 : reciprocal = 16'b0000000000000010;
        15'b000000100010110 : reciprocal = 16'b0000000000000010;
        15'b000000100010111 : reciprocal = 16'b0000000000000010;
        15'b000000100011000 : reciprocal = 16'b0000000000000010;
        15'b000000100011001 : reciprocal = 16'b0000000000000010;
        15'b000000100011010 : reciprocal = 16'b0000000000000010;
        15'b000000100011011 : reciprocal = 16'b0000000000000010;
        15'b000000100011100 : reciprocal = 16'b0000000000000010;
        15'b000000100011101 : reciprocal = 16'b0000000000000010;
        15'b000000100011110 : reciprocal = 16'b0000000000000010;
        15'b000000100011111 : reciprocal = 16'b0000000000000010;
        15'b000000100100000 : reciprocal = 16'b0000000000000010;
        15'b000000100100001 : reciprocal = 16'b0000000000000010;
        15'b000000100100010 : reciprocal = 16'b0000000000000010;
        15'b000000100100011 : reciprocal = 16'b0000000000000010;
        15'b000000100100100 : reciprocal = 16'b0000000000000010;
        15'b000000100100101 : reciprocal = 16'b0000000000000010;
        15'b000000100100110 : reciprocal = 16'b0000000000000010;
        15'b000000100100111 : reciprocal = 16'b0000000000000010;
        15'b000000100101000 : reciprocal = 16'b0000000000000010;
        15'b000000100101001 : reciprocal = 16'b0000000000000010;
        15'b000000100101010 : reciprocal = 16'b0000000000000010;
        15'b000000100101011 : reciprocal = 16'b0000000000000010;
        15'b000000100101100 : reciprocal = 16'b0000000000000010;
        15'b000000100101101 : reciprocal = 16'b0000000000000010;
        15'b000000100101110 : reciprocal = 16'b0000000000000010;
        15'b000000100101111 : reciprocal = 16'b0000000000000010;
        15'b000000100110000 : reciprocal = 16'b0000000000000010;
        15'b000000100110001 : reciprocal = 16'b0000000000000010;
        15'b000000100110010 : reciprocal = 16'b0000000000000010;
        15'b000000100110011 : reciprocal = 16'b0000000000000010;
        15'b000000100110100 : reciprocal = 16'b0000000000000010;
        15'b000000100110101 : reciprocal = 16'b0000000000000010;
        15'b000000100110110 : reciprocal = 16'b0000000000000010;
        15'b000000100110111 : reciprocal = 16'b0000000000000010;
        15'b000000100111000 : reciprocal = 16'b0000000000000010;
        15'b000000100111001 : reciprocal = 16'b0000000000000010;
        15'b000000100111010 : reciprocal = 16'b0000000000000010;
        15'b000000100111011 : reciprocal = 16'b0000000000000010;
        15'b000000100111100 : reciprocal = 16'b0000000000000010;
        15'b000000100111101 : reciprocal = 16'b0000000000000010;
        15'b000000100111110 : reciprocal = 16'b0000000000000010;
        15'b000000100111111 : reciprocal = 16'b0000000000000010;
        15'b000000101000000 : reciprocal = 16'b0000000000000010;
        15'b000000101000001 : reciprocal = 16'b0000000000000010;
        15'b000000101000010 : reciprocal = 16'b0000000000000010;
        15'b000000101000011 : reciprocal = 16'b0000000000000010;
        15'b000000101000100 : reciprocal = 16'b0000000000000010;
        15'b000000101000101 : reciprocal = 16'b0000000000000010;
        15'b000000101000110 : reciprocal = 16'b0000000000000010;
        15'b000000101000111 : reciprocal = 16'b0000000000000010;
        15'b000000101001000 : reciprocal = 16'b0000000000000010;
        15'b000000101001001 : reciprocal = 16'b0000000000000010;
        15'b000000101001010 : reciprocal = 16'b0000000000000010;
        15'b000000101001011 : reciprocal = 16'b0000000000000010;
        15'b000000101001100 : reciprocal = 16'b0000000000000010;
        15'b000000101001101 : reciprocal = 16'b0000000000000010;
        15'b000000101001110 : reciprocal = 16'b0000000000000010;
        15'b000000101001111 : reciprocal = 16'b0000000000000010;
        15'b000000101010000 : reciprocal = 16'b0000000000000010;
        15'b000000101010001 : reciprocal = 16'b0000000000000010;
        15'b000000101010010 : reciprocal = 16'b0000000000000010;
        15'b000000101010011 : reciprocal = 16'b0000000000000010;
        15'b000000101010100 : reciprocal = 16'b0000000000000010;
        15'b000000101010101 : reciprocal = 16'b0000000000000010;
        15'b000000101010110 : reciprocal = 16'b0000000000000001;
        15'b000000101010111 : reciprocal = 16'b0000000000000001;
        15'b000000101011000 : reciprocal = 16'b0000000000000001;
        15'b000000101011001 : reciprocal = 16'b0000000000000001;
        15'b000000101011010 : reciprocal = 16'b0000000000000001;
        15'b000000101011011 : reciprocal = 16'b0000000000000001;
        15'b000000101011100 : reciprocal = 16'b0000000000000001;
        15'b000000101011101 : reciprocal = 16'b0000000000000001;
        15'b000000101011110 : reciprocal = 16'b0000000000000001;
        15'b000000101011111 : reciprocal = 16'b0000000000000001;
        15'b000000101100000 : reciprocal = 16'b0000000000000001;
        15'b000000101100001 : reciprocal = 16'b0000000000000001;
        15'b000000101100010 : reciprocal = 16'b0000000000000001;
        15'b000000101100011 : reciprocal = 16'b0000000000000001;
        15'b000000101100100 : reciprocal = 16'b0000000000000001;
        15'b000000101100101 : reciprocal = 16'b0000000000000001;
        15'b000000101100110 : reciprocal = 16'b0000000000000001;
        15'b000000101100111 : reciprocal = 16'b0000000000000001;
        15'b000000101101000 : reciprocal = 16'b0000000000000001;
        15'b000000101101001 : reciprocal = 16'b0000000000000001;
        15'b000000101101010 : reciprocal = 16'b0000000000000001;
        15'b000000101101011 : reciprocal = 16'b0000000000000001;
        15'b000000101101100 : reciprocal = 16'b0000000000000001;
        15'b000000101101101 : reciprocal = 16'b0000000000000001;
        15'b000000101101110 : reciprocal = 16'b0000000000000001;
        15'b000000101101111 : reciprocal = 16'b0000000000000001;
        15'b000000101110000 : reciprocal = 16'b0000000000000001;
        15'b000000101110001 : reciprocal = 16'b0000000000000001;
        15'b000000101110010 : reciprocal = 16'b0000000000000001;
        15'b000000101110011 : reciprocal = 16'b0000000000000001;
        15'b000000101110100 : reciprocal = 16'b0000000000000001;
        15'b000000101110101 : reciprocal = 16'b0000000000000001;
        15'b000000101110110 : reciprocal = 16'b0000000000000001;
        15'b000000101110111 : reciprocal = 16'b0000000000000001;
        15'b000000101111000 : reciprocal = 16'b0000000000000001;
        15'b000000101111001 : reciprocal = 16'b0000000000000001;
        15'b000000101111010 : reciprocal = 16'b0000000000000001;
        15'b000000101111011 : reciprocal = 16'b0000000000000001;
        15'b000000101111100 : reciprocal = 16'b0000000000000001;
        15'b000000101111101 : reciprocal = 16'b0000000000000001;
        15'b000000101111110 : reciprocal = 16'b0000000000000001;
        15'b000000101111111 : reciprocal = 16'b0000000000000001;
        15'b000000110000000 : reciprocal = 16'b0000000000000001;
        15'b000000110000001 : reciprocal = 16'b0000000000000001;
        15'b000000110000010 : reciprocal = 16'b0000000000000001;
        15'b000000110000011 : reciprocal = 16'b0000000000000001;
        15'b000000110000100 : reciprocal = 16'b0000000000000001;
        15'b000000110000101 : reciprocal = 16'b0000000000000001;
        15'b000000110000110 : reciprocal = 16'b0000000000000001;
        15'b000000110000111 : reciprocal = 16'b0000000000000001;
        15'b000000110001000 : reciprocal = 16'b0000000000000001;
        15'b000000110001001 : reciprocal = 16'b0000000000000001;
        15'b000000110001010 : reciprocal = 16'b0000000000000001;
        15'b000000110001011 : reciprocal = 16'b0000000000000001;
        15'b000000110001100 : reciprocal = 16'b0000000000000001;
        15'b000000110001101 : reciprocal = 16'b0000000000000001;
        15'b000000110001110 : reciprocal = 16'b0000000000000001;
        15'b000000110001111 : reciprocal = 16'b0000000000000001;
        15'b000000110010000 : reciprocal = 16'b0000000000000001;
        15'b000000110010001 : reciprocal = 16'b0000000000000001;
        15'b000000110010010 : reciprocal = 16'b0000000000000001;
        15'b000000110010011 : reciprocal = 16'b0000000000000001;
        15'b000000110010100 : reciprocal = 16'b0000000000000001;
        15'b000000110010101 : reciprocal = 16'b0000000000000001;
        15'b000000110010110 : reciprocal = 16'b0000000000000001;
        15'b000000110010111 : reciprocal = 16'b0000000000000001;
        15'b000000110011000 : reciprocal = 16'b0000000000000001;
        15'b000000110011001 : reciprocal = 16'b0000000000000001;
        15'b000000110011010 : reciprocal = 16'b0000000000000001;
        15'b000000110011011 : reciprocal = 16'b0000000000000001;
        15'b000000110011100 : reciprocal = 16'b0000000000000001;
        15'b000000110011101 : reciprocal = 16'b0000000000000001;
        15'b000000110011110 : reciprocal = 16'b0000000000000001;
        15'b000000110011111 : reciprocal = 16'b0000000000000001;
        15'b000000110100000 : reciprocal = 16'b0000000000000001;
        15'b000000110100001 : reciprocal = 16'b0000000000000001;
        15'b000000110100010 : reciprocal = 16'b0000000000000001;
        15'b000000110100011 : reciprocal = 16'b0000000000000001;
        15'b000000110100100 : reciprocal = 16'b0000000000000001;
        15'b000000110100101 : reciprocal = 16'b0000000000000001;
        15'b000000110100110 : reciprocal = 16'b0000000000000001;
        15'b000000110100111 : reciprocal = 16'b0000000000000001;
        15'b000000110101000 : reciprocal = 16'b0000000000000001;
        15'b000000110101001 : reciprocal = 16'b0000000000000001;
        15'b000000110101010 : reciprocal = 16'b0000000000000001;
        15'b000000110101011 : reciprocal = 16'b0000000000000001;
        15'b000000110101100 : reciprocal = 16'b0000000000000001;
        15'b000000110101101 : reciprocal = 16'b0000000000000001;
        15'b000000110101110 : reciprocal = 16'b0000000000000001;
        15'b000000110101111 : reciprocal = 16'b0000000000000001;
        15'b000000110110000 : reciprocal = 16'b0000000000000001;
        15'b000000110110001 : reciprocal = 16'b0000000000000001;
        15'b000000110110010 : reciprocal = 16'b0000000000000001;
        15'b000000110110011 : reciprocal = 16'b0000000000000001;
        15'b000000110110100 : reciprocal = 16'b0000000000000001;
        15'b000000110110101 : reciprocal = 16'b0000000000000001;
        15'b000000110110110 : reciprocal = 16'b0000000000000001;
        15'b000000110110111 : reciprocal = 16'b0000000000000001;
        15'b000000110111000 : reciprocal = 16'b0000000000000001;
        15'b000000110111001 : reciprocal = 16'b0000000000000001;
        15'b000000110111010 : reciprocal = 16'b0000000000000001;
        15'b000000110111011 : reciprocal = 16'b0000000000000001;
        15'b000000110111100 : reciprocal = 16'b0000000000000001;
        15'b000000110111101 : reciprocal = 16'b0000000000000001;
        15'b000000110111110 : reciprocal = 16'b0000000000000001;
        15'b000000110111111 : reciprocal = 16'b0000000000000001;
        15'b000000111000000 : reciprocal = 16'b0000000000000001;
        15'b000000111000001 : reciprocal = 16'b0000000000000001;
        15'b000000111000010 : reciprocal = 16'b0000000000000001;
        15'b000000111000011 : reciprocal = 16'b0000000000000001;
        15'b000000111000100 : reciprocal = 16'b0000000000000001;
        15'b000000111000101 : reciprocal = 16'b0000000000000001;
        15'b000000111000110 : reciprocal = 16'b0000000000000001;
        15'b000000111000111 : reciprocal = 16'b0000000000000001;
        15'b000000111001000 : reciprocal = 16'b0000000000000001;
        15'b000000111001001 : reciprocal = 16'b0000000000000001;
        15'b000000111001010 : reciprocal = 16'b0000000000000001;
        15'b000000111001011 : reciprocal = 16'b0000000000000001;
        15'b000000111001100 : reciprocal = 16'b0000000000000001;
        15'b000000111001101 : reciprocal = 16'b0000000000000001;
        15'b000000111001110 : reciprocal = 16'b0000000000000001;
        15'b000000111001111 : reciprocal = 16'b0000000000000001;
        15'b000000111010000 : reciprocal = 16'b0000000000000001;
        15'b000000111010001 : reciprocal = 16'b0000000000000001;
        15'b000000111010010 : reciprocal = 16'b0000000000000001;
        15'b000000111010011 : reciprocal = 16'b0000000000000001;
        15'b000000111010100 : reciprocal = 16'b0000000000000001;
        15'b000000111010101 : reciprocal = 16'b0000000000000001;
        15'b000000111010110 : reciprocal = 16'b0000000000000001;
        15'b000000111010111 : reciprocal = 16'b0000000000000001;
        15'b000000111011000 : reciprocal = 16'b0000000000000001;
        15'b000000111011001 : reciprocal = 16'b0000000000000001;
        15'b000000111011010 : reciprocal = 16'b0000000000000001;
        15'b000000111011011 : reciprocal = 16'b0000000000000001;
        15'b000000111011100 : reciprocal = 16'b0000000000000001;
        15'b000000111011101 : reciprocal = 16'b0000000000000001;
        15'b000000111011110 : reciprocal = 16'b0000000000000001;
        15'b000000111011111 : reciprocal = 16'b0000000000000001;
        15'b000000111100000 : reciprocal = 16'b0000000000000001;
        15'b000000111100001 : reciprocal = 16'b0000000000000001;
        15'b000000111100010 : reciprocal = 16'b0000000000000001;
        15'b000000111100011 : reciprocal = 16'b0000000000000001;
        15'b000000111100100 : reciprocal = 16'b0000000000000001;
        15'b000000111100101 : reciprocal = 16'b0000000000000001;
        15'b000000111100110 : reciprocal = 16'b0000000000000001;
        15'b000000111100111 : reciprocal = 16'b0000000000000001;
        15'b000000111101000 : reciprocal = 16'b0000000000000001;
        15'b000000111101001 : reciprocal = 16'b0000000000000001;
        15'b000000111101010 : reciprocal = 16'b0000000000000001;
        15'b000000111101011 : reciprocal = 16'b0000000000000001;
        15'b000000111101100 : reciprocal = 16'b0000000000000001;
        15'b000000111101101 : reciprocal = 16'b0000000000000001;
        15'b000000111101110 : reciprocal = 16'b0000000000000001;
        15'b000000111101111 : reciprocal = 16'b0000000000000001;
        15'b000000111110000 : reciprocal = 16'b0000000000000001;
        15'b000000111110001 : reciprocal = 16'b0000000000000001;
        15'b000000111110010 : reciprocal = 16'b0000000000000001;
        15'b000000111110011 : reciprocal = 16'b0000000000000001;
        15'b000000111110100 : reciprocal = 16'b0000000000000001;
        15'b000000111110101 : reciprocal = 16'b0000000000000001;
        15'b000000111110110 : reciprocal = 16'b0000000000000001;
        15'b000000111110111 : reciprocal = 16'b0000000000000001;
        15'b000000111111000 : reciprocal = 16'b0000000000000001;
        15'b000000111111001 : reciprocal = 16'b0000000000000001;
        15'b000000111111010 : reciprocal = 16'b0000000000000001;
        15'b000000111111011 : reciprocal = 16'b0000000000000001;
        15'b000000111111100 : reciprocal = 16'b0000000000000001;
        15'b000000111111101 : reciprocal = 16'b0000000000000001;
        15'b000000111111110 : reciprocal = 16'b0000000000000001;
        15'b000000111111111 : reciprocal = 16'b0000000000000001;
        15'b000001000000000 : reciprocal = 16'b0000000000000001;
        15'b000001000000001 : reciprocal = 16'b0000000000000001;
        15'b000001000000010 : reciprocal = 16'b0000000000000001;
        15'b000001000000011 : reciprocal = 16'b0000000000000001;
        15'b000001000000100 : reciprocal = 16'b0000000000000001;
        15'b000001000000101 : reciprocal = 16'b0000000000000001;
        15'b000001000000110 : reciprocal = 16'b0000000000000001;
        15'b000001000000111 : reciprocal = 16'b0000000000000001;
        15'b000001000001000 : reciprocal = 16'b0000000000000001;
        15'b000001000001001 : reciprocal = 16'b0000000000000001;
        15'b000001000001010 : reciprocal = 16'b0000000000000001;
        15'b000001000001011 : reciprocal = 16'b0000000000000001;
        15'b000001000001100 : reciprocal = 16'b0000000000000001;
        15'b000001000001101 : reciprocal = 16'b0000000000000001;
        15'b000001000001110 : reciprocal = 16'b0000000000000001;
        15'b000001000001111 : reciprocal = 16'b0000000000000001;
        15'b000001000010000 : reciprocal = 16'b0000000000000001;
        15'b000001000010001 : reciprocal = 16'b0000000000000001;
        15'b000001000010010 : reciprocal = 16'b0000000000000001;
        15'b000001000010011 : reciprocal = 16'b0000000000000001;
        15'b000001000010100 : reciprocal = 16'b0000000000000001;
        15'b000001000010101 : reciprocal = 16'b0000000000000001;
        15'b000001000010110 : reciprocal = 16'b0000000000000001;
        15'b000001000010111 : reciprocal = 16'b0000000000000001;
        15'b000001000011000 : reciprocal = 16'b0000000000000001;
        15'b000001000011001 : reciprocal = 16'b0000000000000001;
        15'b000001000011010 : reciprocal = 16'b0000000000000001;
        15'b000001000011011 : reciprocal = 16'b0000000000000001;
        15'b000001000011100 : reciprocal = 16'b0000000000000001;
        15'b000001000011101 : reciprocal = 16'b0000000000000001;
        15'b000001000011110 : reciprocal = 16'b0000000000000001;
        15'b000001000011111 : reciprocal = 16'b0000000000000001;
        15'b000001000100000 : reciprocal = 16'b0000000000000001;
        15'b000001000100001 : reciprocal = 16'b0000000000000001;
        15'b000001000100010 : reciprocal = 16'b0000000000000001;
        15'b000001000100011 : reciprocal = 16'b0000000000000001;
        15'b000001000100100 : reciprocal = 16'b0000000000000001;
        15'b000001000100101 : reciprocal = 16'b0000000000000001;
        15'b000001000100110 : reciprocal = 16'b0000000000000001;
        15'b000001000100111 : reciprocal = 16'b0000000000000001;
        15'b000001000101000 : reciprocal = 16'b0000000000000001;
        15'b000001000101001 : reciprocal = 16'b0000000000000001;
        15'b000001000101010 : reciprocal = 16'b0000000000000001;
        15'b000001000101011 : reciprocal = 16'b0000000000000001;
        15'b000001000101100 : reciprocal = 16'b0000000000000001;
        15'b000001000101101 : reciprocal = 16'b0000000000000001;
        15'b000001000101110 : reciprocal = 16'b0000000000000001;
        15'b000001000101111 : reciprocal = 16'b0000000000000001;
        15'b000001000110000 : reciprocal = 16'b0000000000000001;
        15'b000001000110001 : reciprocal = 16'b0000000000000001;
        15'b000001000110010 : reciprocal = 16'b0000000000000001;
        15'b000001000110011 : reciprocal = 16'b0000000000000001;
        15'b000001000110100 : reciprocal = 16'b0000000000000001;
        15'b000001000110101 : reciprocal = 16'b0000000000000001;
        15'b000001000110110 : reciprocal = 16'b0000000000000001;
        15'b000001000110111 : reciprocal = 16'b0000000000000001;
        15'b000001000111000 : reciprocal = 16'b0000000000000001;
        15'b000001000111001 : reciprocal = 16'b0000000000000001;
        15'b000001000111010 : reciprocal = 16'b0000000000000001;
        15'b000001000111011 : reciprocal = 16'b0000000000000001;
        15'b000001000111100 : reciprocal = 16'b0000000000000001;
        15'b000001000111101 : reciprocal = 16'b0000000000000001;
        15'b000001000111110 : reciprocal = 16'b0000000000000001;
        15'b000001000111111 : reciprocal = 16'b0000000000000001;
        15'b000001001000000 : reciprocal = 16'b0000000000000001;
        15'b000001001000001 : reciprocal = 16'b0000000000000001;
        15'b000001001000010 : reciprocal = 16'b0000000000000001;
        15'b000001001000011 : reciprocal = 16'b0000000000000001;
        15'b000001001000100 : reciprocal = 16'b0000000000000001;
        15'b000001001000101 : reciprocal = 16'b0000000000000001;
        15'b000001001000110 : reciprocal = 16'b0000000000000001;
        15'b000001001000111 : reciprocal = 16'b0000000000000001;
        15'b000001001001000 : reciprocal = 16'b0000000000000001;
        15'b000001001001001 : reciprocal = 16'b0000000000000001;
        15'b000001001001010 : reciprocal = 16'b0000000000000001;
        15'b000001001001011 : reciprocal = 16'b0000000000000001;
        15'b000001001001100 : reciprocal = 16'b0000000000000001;
        15'b000001001001101 : reciprocal = 16'b0000000000000001;
        15'b000001001001110 : reciprocal = 16'b0000000000000001;
        15'b000001001001111 : reciprocal = 16'b0000000000000001;
        15'b000001001010000 : reciprocal = 16'b0000000000000001;
        15'b000001001010001 : reciprocal = 16'b0000000000000001;
        15'b000001001010010 : reciprocal = 16'b0000000000000001;
        15'b000001001010011 : reciprocal = 16'b0000000000000001;
        15'b000001001010100 : reciprocal = 16'b0000000000000001;
        15'b000001001010101 : reciprocal = 16'b0000000000000001;
        15'b000001001010110 : reciprocal = 16'b0000000000000001;
        15'b000001001010111 : reciprocal = 16'b0000000000000001;
        15'b000001001011000 : reciprocal = 16'b0000000000000001;
        15'b000001001011001 : reciprocal = 16'b0000000000000001;
        15'b000001001011010 : reciprocal = 16'b0000000000000001;
        15'b000001001011011 : reciprocal = 16'b0000000000000001;
        15'b000001001011100 : reciprocal = 16'b0000000000000001;
        15'b000001001011101 : reciprocal = 16'b0000000000000001;
        15'b000001001011110 : reciprocal = 16'b0000000000000001;
        15'b000001001011111 : reciprocal = 16'b0000000000000001;
        15'b000001001100000 : reciprocal = 16'b0000000000000001;
        15'b000001001100001 : reciprocal = 16'b0000000000000001;
        15'b000001001100010 : reciprocal = 16'b0000000000000001;
        15'b000001001100011 : reciprocal = 16'b0000000000000001;
        15'b000001001100100 : reciprocal = 16'b0000000000000001;
        15'b000001001100101 : reciprocal = 16'b0000000000000001;
        15'b000001001100110 : reciprocal = 16'b0000000000000001;
        15'b000001001100111 : reciprocal = 16'b0000000000000001;
        15'b000001001101000 : reciprocal = 16'b0000000000000001;
        15'b000001001101001 : reciprocal = 16'b0000000000000001;
        15'b000001001101010 : reciprocal = 16'b0000000000000001;
        15'b000001001101011 : reciprocal = 16'b0000000000000001;
        15'b000001001101100 : reciprocal = 16'b0000000000000001;
        15'b000001001101101 : reciprocal = 16'b0000000000000001;
        15'b000001001101110 : reciprocal = 16'b0000000000000001;
        15'b000001001101111 : reciprocal = 16'b0000000000000001;
        15'b000001001110000 : reciprocal = 16'b0000000000000001;
        15'b000001001110001 : reciprocal = 16'b0000000000000001;
        15'b000001001110010 : reciprocal = 16'b0000000000000001;
        15'b000001001110011 : reciprocal = 16'b0000000000000001;
        15'b000001001110100 : reciprocal = 16'b0000000000000001;
        15'b000001001110101 : reciprocal = 16'b0000000000000001;
        15'b000001001110110 : reciprocal = 16'b0000000000000001;
        15'b000001001110111 : reciprocal = 16'b0000000000000001;
        15'b000001001111000 : reciprocal = 16'b0000000000000001;
        15'b000001001111001 : reciprocal = 16'b0000000000000001;
        15'b000001001111010 : reciprocal = 16'b0000000000000001;
        15'b000001001111011 : reciprocal = 16'b0000000000000001;
        15'b000001001111100 : reciprocal = 16'b0000000000000001;
        15'b000001001111101 : reciprocal = 16'b0000000000000001;
        15'b000001001111110 : reciprocal = 16'b0000000000000001;
        15'b000001001111111 : reciprocal = 16'b0000000000000001;
        15'b000001010000000 : reciprocal = 16'b0000000000000001;
        15'b000001010000001 : reciprocal = 16'b0000000000000001;
        15'b000001010000010 : reciprocal = 16'b0000000000000001;
        15'b000001010000011 : reciprocal = 16'b0000000000000001;
        15'b000001010000100 : reciprocal = 16'b0000000000000001;
        15'b000001010000101 : reciprocal = 16'b0000000000000001;
        15'b000001010000110 : reciprocal = 16'b0000000000000001;
        15'b000001010000111 : reciprocal = 16'b0000000000000001;
        15'b000001010001000 : reciprocal = 16'b0000000000000001;
        15'b000001010001001 : reciprocal = 16'b0000000000000001;
        15'b000001010001010 : reciprocal = 16'b0000000000000001;
        15'b000001010001011 : reciprocal = 16'b0000000000000001;
        15'b000001010001100 : reciprocal = 16'b0000000000000001;
        15'b000001010001101 : reciprocal = 16'b0000000000000001;
        15'b000001010001110 : reciprocal = 16'b0000000000000001;
        15'b000001010001111 : reciprocal = 16'b0000000000000001;
        15'b000001010010000 : reciprocal = 16'b0000000000000001;
        15'b000001010010001 : reciprocal = 16'b0000000000000001;
        15'b000001010010010 : reciprocal = 16'b0000000000000001;
        15'b000001010010011 : reciprocal = 16'b0000000000000001;
        15'b000001010010100 : reciprocal = 16'b0000000000000001;
        15'b000001010010101 : reciprocal = 16'b0000000000000001;
        15'b000001010010110 : reciprocal = 16'b0000000000000001;
        15'b000001010010111 : reciprocal = 16'b0000000000000001;
        15'b000001010011000 : reciprocal = 16'b0000000000000001;
        15'b000001010011001 : reciprocal = 16'b0000000000000001;
        15'b000001010011010 : reciprocal = 16'b0000000000000001;
        15'b000001010011011 : reciprocal = 16'b0000000000000001;
        15'b000001010011100 : reciprocal = 16'b0000000000000001;
        15'b000001010011101 : reciprocal = 16'b0000000000000001;
        15'b000001010011110 : reciprocal = 16'b0000000000000001;
        15'b000001010011111 : reciprocal = 16'b0000000000000001;
        15'b000001010100000 : reciprocal = 16'b0000000000000001;
        15'b000001010100001 : reciprocal = 16'b0000000000000001;
        15'b000001010100010 : reciprocal = 16'b0000000000000001;
        15'b000001010100011 : reciprocal = 16'b0000000000000001;
        15'b000001010100100 : reciprocal = 16'b0000000000000001;
        15'b000001010100101 : reciprocal = 16'b0000000000000001;
        15'b000001010100110 : reciprocal = 16'b0000000000000001;
        15'b000001010100111 : reciprocal = 16'b0000000000000001;
        15'b000001010101000 : reciprocal = 16'b0000000000000001;
        15'b000001010101001 : reciprocal = 16'b0000000000000001;
        15'b000001010101010 : reciprocal = 16'b0000000000000001;
        15'b000001010101011 : reciprocal = 16'b0000000000000001;
        15'b000001010101100 : reciprocal = 16'b0000000000000001;
        15'b000001010101101 : reciprocal = 16'b0000000000000001;
        15'b000001010101110 : reciprocal = 16'b0000000000000001;
        15'b000001010101111 : reciprocal = 16'b0000000000000001;
        15'b000001010110000 : reciprocal = 16'b0000000000000001;
        15'b000001010110001 : reciprocal = 16'b0000000000000001;
        15'b000001010110010 : reciprocal = 16'b0000000000000001;
        15'b000001010110011 : reciprocal = 16'b0000000000000001;
        15'b000001010110100 : reciprocal = 16'b0000000000000001;
        15'b000001010110101 : reciprocal = 16'b0000000000000001;
        15'b000001010110110 : reciprocal = 16'b0000000000000001;
        15'b000001010110111 : reciprocal = 16'b0000000000000001;
        15'b000001010111000 : reciprocal = 16'b0000000000000001;
        15'b000001010111001 : reciprocal = 16'b0000000000000001;
        15'b000001010111010 : reciprocal = 16'b0000000000000001;
        15'b000001010111011 : reciprocal = 16'b0000000000000001;
        15'b000001010111100 : reciprocal = 16'b0000000000000001;
        15'b000001010111101 : reciprocal = 16'b0000000000000001;
        15'b000001010111110 : reciprocal = 16'b0000000000000001;
        15'b000001010111111 : reciprocal = 16'b0000000000000001;
        15'b000001011000000 : reciprocal = 16'b0000000000000001;
        15'b000001011000001 : reciprocal = 16'b0000000000000001;
        15'b000001011000010 : reciprocal = 16'b0000000000000001;
        15'b000001011000011 : reciprocal = 16'b0000000000000001;
        15'b000001011000100 : reciprocal = 16'b0000000000000001;
        15'b000001011000101 : reciprocal = 16'b0000000000000001;
        15'b000001011000110 : reciprocal = 16'b0000000000000001;
        15'b000001011000111 : reciprocal = 16'b0000000000000001;
        15'b000001011001000 : reciprocal = 16'b0000000000000001;
        15'b000001011001001 : reciprocal = 16'b0000000000000001;
        15'b000001011001010 : reciprocal = 16'b0000000000000001;
        15'b000001011001011 : reciprocal = 16'b0000000000000001;
        15'b000001011001100 : reciprocal = 16'b0000000000000001;
        15'b000001011001101 : reciprocal = 16'b0000000000000001;
        15'b000001011001110 : reciprocal = 16'b0000000000000001;
        15'b000001011001111 : reciprocal = 16'b0000000000000001;
        15'b000001011010000 : reciprocal = 16'b0000000000000001;
        15'b000001011010001 : reciprocal = 16'b0000000000000001;
        15'b000001011010010 : reciprocal = 16'b0000000000000001;
        15'b000001011010011 : reciprocal = 16'b0000000000000001;
        15'b000001011010100 : reciprocal = 16'b0000000000000001;
        15'b000001011010101 : reciprocal = 16'b0000000000000001;
        15'b000001011010110 : reciprocal = 16'b0000000000000001;
        15'b000001011010111 : reciprocal = 16'b0000000000000001;
        15'b000001011011000 : reciprocal = 16'b0000000000000001;
        15'b000001011011001 : reciprocal = 16'b0000000000000001;
        15'b000001011011010 : reciprocal = 16'b0000000000000001;
        15'b000001011011011 : reciprocal = 16'b0000000000000001;
        15'b000001011011100 : reciprocal = 16'b0000000000000001;
        15'b000001011011101 : reciprocal = 16'b0000000000000001;
        15'b000001011011110 : reciprocal = 16'b0000000000000001;
        15'b000001011011111 : reciprocal = 16'b0000000000000001;
        15'b000001011100000 : reciprocal = 16'b0000000000000001;
        15'b000001011100001 : reciprocal = 16'b0000000000000001;
        15'b000001011100010 : reciprocal = 16'b0000000000000001;
        15'b000001011100011 : reciprocal = 16'b0000000000000001;
        15'b000001011100100 : reciprocal = 16'b0000000000000001;
        15'b000001011100101 : reciprocal = 16'b0000000000000001;
        15'b000001011100110 : reciprocal = 16'b0000000000000001;
        15'b000001011100111 : reciprocal = 16'b0000000000000001;
        15'b000001011101000 : reciprocal = 16'b0000000000000001;
        15'b000001011101001 : reciprocal = 16'b0000000000000001;
        15'b000001011101010 : reciprocal = 16'b0000000000000001;
        15'b000001011101011 : reciprocal = 16'b0000000000000001;
        15'b000001011101100 : reciprocal = 16'b0000000000000001;
        15'b000001011101101 : reciprocal = 16'b0000000000000001;
        15'b000001011101110 : reciprocal = 16'b0000000000000001;
        15'b000001011101111 : reciprocal = 16'b0000000000000001;
        15'b000001011110000 : reciprocal = 16'b0000000000000001;
        15'b000001011110001 : reciprocal = 16'b0000000000000001;
        15'b000001011110010 : reciprocal = 16'b0000000000000001;
        15'b000001011110011 : reciprocal = 16'b0000000000000001;
        15'b000001011110100 : reciprocal = 16'b0000000000000001;
        15'b000001011110101 : reciprocal = 16'b0000000000000001;
        15'b000001011110110 : reciprocal = 16'b0000000000000001;
        15'b000001011110111 : reciprocal = 16'b0000000000000001;
        15'b000001011111000 : reciprocal = 16'b0000000000000001;
        15'b000001011111001 : reciprocal = 16'b0000000000000001;
        15'b000001011111010 : reciprocal = 16'b0000000000000001;
        15'b000001011111011 : reciprocal = 16'b0000000000000001;
        15'b000001011111100 : reciprocal = 16'b0000000000000001;
        15'b000001011111101 : reciprocal = 16'b0000000000000001;
        15'b000001011111110 : reciprocal = 16'b0000000000000001;
        15'b000001011111111 : reciprocal = 16'b0000000000000001;
        15'b000001100000000 : reciprocal = 16'b0000000000000001;
        15'b000001100000001 : reciprocal = 16'b0000000000000001;
        15'b000001100000010 : reciprocal = 16'b0000000000000001;
        15'b000001100000011 : reciprocal = 16'b0000000000000001;
        15'b000001100000100 : reciprocal = 16'b0000000000000001;
        15'b000001100000101 : reciprocal = 16'b0000000000000001;
        15'b000001100000110 : reciprocal = 16'b0000000000000001;
        15'b000001100000111 : reciprocal = 16'b0000000000000001;
        15'b000001100001000 : reciprocal = 16'b0000000000000001;
        15'b000001100001001 : reciprocal = 16'b0000000000000001;
        15'b000001100001010 : reciprocal = 16'b0000000000000001;
        15'b000001100001011 : reciprocal = 16'b0000000000000001;
        15'b000001100001100 : reciprocal = 16'b0000000000000001;
        15'b000001100001101 : reciprocal = 16'b0000000000000001;
        15'b000001100001110 : reciprocal = 16'b0000000000000001;
        15'b000001100001111 : reciprocal = 16'b0000000000000001;
        15'b000001100010000 : reciprocal = 16'b0000000000000001;
        15'b000001100010001 : reciprocal = 16'b0000000000000001;
        15'b000001100010010 : reciprocal = 16'b0000000000000001;
        15'b000001100010011 : reciprocal = 16'b0000000000000001;
        15'b000001100010100 : reciprocal = 16'b0000000000000001;
        15'b000001100010101 : reciprocal = 16'b0000000000000001;
        15'b000001100010110 : reciprocal = 16'b0000000000000001;
        15'b000001100010111 : reciprocal = 16'b0000000000000001;
        15'b000001100011000 : reciprocal = 16'b0000000000000001;
        15'b000001100011001 : reciprocal = 16'b0000000000000001;
        15'b000001100011010 : reciprocal = 16'b0000000000000001;
        15'b000001100011011 : reciprocal = 16'b0000000000000001;
        15'b000001100011100 : reciprocal = 16'b0000000000000001;
        15'b000001100011101 : reciprocal = 16'b0000000000000001;
        15'b000001100011110 : reciprocal = 16'b0000000000000001;
        15'b000001100011111 : reciprocal = 16'b0000000000000001;
        15'b000001100100000 : reciprocal = 16'b0000000000000001;
        15'b000001100100001 : reciprocal = 16'b0000000000000001;
        15'b000001100100010 : reciprocal = 16'b0000000000000001;
        15'b000001100100011 : reciprocal = 16'b0000000000000001;
        15'b000001100100100 : reciprocal = 16'b0000000000000001;
        15'b000001100100101 : reciprocal = 16'b0000000000000001;
        15'b000001100100110 : reciprocal = 16'b0000000000000001;
        15'b000001100100111 : reciprocal = 16'b0000000000000001;
        15'b000001100101000 : reciprocal = 16'b0000000000000001;
        15'b000001100101001 : reciprocal = 16'b0000000000000001;
        15'b000001100101010 : reciprocal = 16'b0000000000000001;
        15'b000001100101011 : reciprocal = 16'b0000000000000001;
        15'b000001100101100 : reciprocal = 16'b0000000000000001;
        15'b000001100101101 : reciprocal = 16'b0000000000000001;
        15'b000001100101110 : reciprocal = 16'b0000000000000001;
        15'b000001100101111 : reciprocal = 16'b0000000000000001;
        15'b000001100110000 : reciprocal = 16'b0000000000000001;
        15'b000001100110001 : reciprocal = 16'b0000000000000001;
        15'b000001100110010 : reciprocal = 16'b0000000000000001;
        15'b000001100110011 : reciprocal = 16'b0000000000000001;
        15'b000001100110100 : reciprocal = 16'b0000000000000001;
        15'b000001100110101 : reciprocal = 16'b0000000000000001;
        15'b000001100110110 : reciprocal = 16'b0000000000000001;
        15'b000001100110111 : reciprocal = 16'b0000000000000001;
        15'b000001100111000 : reciprocal = 16'b0000000000000001;
        15'b000001100111001 : reciprocal = 16'b0000000000000001;
        15'b000001100111010 : reciprocal = 16'b0000000000000001;
        15'b000001100111011 : reciprocal = 16'b0000000000000001;
        15'b000001100111100 : reciprocal = 16'b0000000000000001;
        15'b000001100111101 : reciprocal = 16'b0000000000000001;
        15'b000001100111110 : reciprocal = 16'b0000000000000001;
        15'b000001100111111 : reciprocal = 16'b0000000000000001;
        15'b000001101000000 : reciprocal = 16'b0000000000000001;
        15'b000001101000001 : reciprocal = 16'b0000000000000001;
        15'b000001101000010 : reciprocal = 16'b0000000000000001;
        15'b000001101000011 : reciprocal = 16'b0000000000000001;
        15'b000001101000100 : reciprocal = 16'b0000000000000001;
        15'b000001101000101 : reciprocal = 16'b0000000000000001;
        15'b000001101000110 : reciprocal = 16'b0000000000000001;
        15'b000001101000111 : reciprocal = 16'b0000000000000001;
        15'b000001101001000 : reciprocal = 16'b0000000000000001;
        15'b000001101001001 : reciprocal = 16'b0000000000000001;
        15'b000001101001010 : reciprocal = 16'b0000000000000001;
        15'b000001101001011 : reciprocal = 16'b0000000000000001;
        15'b000001101001100 : reciprocal = 16'b0000000000000001;
        15'b000001101001101 : reciprocal = 16'b0000000000000001;
        15'b000001101001110 : reciprocal = 16'b0000000000000001;
        15'b000001101001111 : reciprocal = 16'b0000000000000001;
        15'b000001101010000 : reciprocal = 16'b0000000000000001;
        15'b000001101010001 : reciprocal = 16'b0000000000000001;
        15'b000001101010010 : reciprocal = 16'b0000000000000001;
        15'b000001101010011 : reciprocal = 16'b0000000000000001;
        15'b000001101010100 : reciprocal = 16'b0000000000000001;
        15'b000001101010101 : reciprocal = 16'b0000000000000001;
        15'b000001101010110 : reciprocal = 16'b0000000000000001;
        15'b000001101010111 : reciprocal = 16'b0000000000000001;
        15'b000001101011000 : reciprocal = 16'b0000000000000001;
        15'b000001101011001 : reciprocal = 16'b0000000000000001;
        15'b000001101011010 : reciprocal = 16'b0000000000000001;
        15'b000001101011011 : reciprocal = 16'b0000000000000001;
        15'b000001101011100 : reciprocal = 16'b0000000000000001;
        15'b000001101011101 : reciprocal = 16'b0000000000000001;
        15'b000001101011110 : reciprocal = 16'b0000000000000001;
        15'b000001101011111 : reciprocal = 16'b0000000000000001;
        15'b000001101100000 : reciprocal = 16'b0000000000000001;
        15'b000001101100001 : reciprocal = 16'b0000000000000001;
        15'b000001101100010 : reciprocal = 16'b0000000000000001;
        15'b000001101100011 : reciprocal = 16'b0000000000000001;
        15'b000001101100100 : reciprocal = 16'b0000000000000001;
        15'b000001101100101 : reciprocal = 16'b0000000000000001;
        15'b000001101100110 : reciprocal = 16'b0000000000000001;
        15'b000001101100111 : reciprocal = 16'b0000000000000001;
        15'b000001101101000 : reciprocal = 16'b0000000000000001;
        15'b000001101101001 : reciprocal = 16'b0000000000000001;
        15'b000001101101010 : reciprocal = 16'b0000000000000001;
        15'b000001101101011 : reciprocal = 16'b0000000000000001;
        15'b000001101101100 : reciprocal = 16'b0000000000000001;
        15'b000001101101101 : reciprocal = 16'b0000000000000001;
        15'b000001101101110 : reciprocal = 16'b0000000000000001;
        15'b000001101101111 : reciprocal = 16'b0000000000000001;
        15'b000001101110000 : reciprocal = 16'b0000000000000001;
        15'b000001101110001 : reciprocal = 16'b0000000000000001;
        15'b000001101110010 : reciprocal = 16'b0000000000000001;
        15'b000001101110011 : reciprocal = 16'b0000000000000001;
        15'b000001101110100 : reciprocal = 16'b0000000000000001;
        15'b000001101110101 : reciprocal = 16'b0000000000000001;
        15'b000001101110110 : reciprocal = 16'b0000000000000001;
        15'b000001101110111 : reciprocal = 16'b0000000000000001;
        15'b000001101111000 : reciprocal = 16'b0000000000000001;
        15'b000001101111001 : reciprocal = 16'b0000000000000001;
        15'b000001101111010 : reciprocal = 16'b0000000000000001;
        15'b000001101111011 : reciprocal = 16'b0000000000000001;
        15'b000001101111100 : reciprocal = 16'b0000000000000001;
        15'b000001101111101 : reciprocal = 16'b0000000000000001;
        15'b000001101111110 : reciprocal = 16'b0000000000000001;
        15'b000001101111111 : reciprocal = 16'b0000000000000001;
        15'b000001110000000 : reciprocal = 16'b0000000000000001;
        15'b000001110000001 : reciprocal = 16'b0000000000000001;
        15'b000001110000010 : reciprocal = 16'b0000000000000001;
        15'b000001110000011 : reciprocal = 16'b0000000000000001;
        15'b000001110000100 : reciprocal = 16'b0000000000000001;
        15'b000001110000101 : reciprocal = 16'b0000000000000001;
        15'b000001110000110 : reciprocal = 16'b0000000000000001;
        15'b000001110000111 : reciprocal = 16'b0000000000000001;
        15'b000001110001000 : reciprocal = 16'b0000000000000001;
        15'b000001110001001 : reciprocal = 16'b0000000000000001;
        15'b000001110001010 : reciprocal = 16'b0000000000000001;
        15'b000001110001011 : reciprocal = 16'b0000000000000001;
        15'b000001110001100 : reciprocal = 16'b0000000000000001;
        15'b000001110001101 : reciprocal = 16'b0000000000000001;
        15'b000001110001110 : reciprocal = 16'b0000000000000001;
        15'b000001110001111 : reciprocal = 16'b0000000000000001;
        15'b000001110010000 : reciprocal = 16'b0000000000000001;
        15'b000001110010001 : reciprocal = 16'b0000000000000001;
        15'b000001110010010 : reciprocal = 16'b0000000000000001;
        15'b000001110010011 : reciprocal = 16'b0000000000000001;
        15'b000001110010100 : reciprocal = 16'b0000000000000001;
        15'b000001110010101 : reciprocal = 16'b0000000000000001;
        15'b000001110010110 : reciprocal = 16'b0000000000000001;
        15'b000001110010111 : reciprocal = 16'b0000000000000001;
        15'b000001110011000 : reciprocal = 16'b0000000000000001;
        15'b000001110011001 : reciprocal = 16'b0000000000000001;
        15'b000001110011010 : reciprocal = 16'b0000000000000001;
        15'b000001110011011 : reciprocal = 16'b0000000000000001;
        15'b000001110011100 : reciprocal = 16'b0000000000000001;
        15'b000001110011101 : reciprocal = 16'b0000000000000001;
        15'b000001110011110 : reciprocal = 16'b0000000000000001;
        15'b000001110011111 : reciprocal = 16'b0000000000000001;
        15'b000001110100000 : reciprocal = 16'b0000000000000001;
        15'b000001110100001 : reciprocal = 16'b0000000000000001;
        15'b000001110100010 : reciprocal = 16'b0000000000000001;
        15'b000001110100011 : reciprocal = 16'b0000000000000001;
        15'b000001110100100 : reciprocal = 16'b0000000000000001;
        15'b000001110100101 : reciprocal = 16'b0000000000000001;
        15'b000001110100110 : reciprocal = 16'b0000000000000001;
        15'b000001110100111 : reciprocal = 16'b0000000000000001;
        15'b000001110101000 : reciprocal = 16'b0000000000000001;
        15'b000001110101001 : reciprocal = 16'b0000000000000001;
        15'b000001110101010 : reciprocal = 16'b0000000000000001;
        15'b000001110101011 : reciprocal = 16'b0000000000000001;
        15'b000001110101100 : reciprocal = 16'b0000000000000001;
        15'b000001110101101 : reciprocal = 16'b0000000000000001;
        15'b000001110101110 : reciprocal = 16'b0000000000000001;
        15'b000001110101111 : reciprocal = 16'b0000000000000001;
        15'b000001110110000 : reciprocal = 16'b0000000000000001;
        15'b000001110110001 : reciprocal = 16'b0000000000000001;
        15'b000001110110010 : reciprocal = 16'b0000000000000001;
        15'b000001110110011 : reciprocal = 16'b0000000000000001;
        15'b000001110110100 : reciprocal = 16'b0000000000000001;
        15'b000001110110101 : reciprocal = 16'b0000000000000001;
        15'b000001110110110 : reciprocal = 16'b0000000000000001;
        15'b000001110110111 : reciprocal = 16'b0000000000000001;
        15'b000001110111000 : reciprocal = 16'b0000000000000001;
        15'b000001110111001 : reciprocal = 16'b0000000000000001;
        15'b000001110111010 : reciprocal = 16'b0000000000000001;
        15'b000001110111011 : reciprocal = 16'b0000000000000001;
        15'b000001110111100 : reciprocal = 16'b0000000000000001;
        15'b000001110111101 : reciprocal = 16'b0000000000000001;
        15'b000001110111110 : reciprocal = 16'b0000000000000001;
        15'b000001110111111 : reciprocal = 16'b0000000000000001;
        15'b000001111000000 : reciprocal = 16'b0000000000000001;
        15'b000001111000001 : reciprocal = 16'b0000000000000001;
        15'b000001111000010 : reciprocal = 16'b0000000000000001;
        15'b000001111000011 : reciprocal = 16'b0000000000000001;
        15'b000001111000100 : reciprocal = 16'b0000000000000001;
        15'b000001111000101 : reciprocal = 16'b0000000000000001;
        15'b000001111000110 : reciprocal = 16'b0000000000000001;
        15'b000001111000111 : reciprocal = 16'b0000000000000001;
        15'b000001111001000 : reciprocal = 16'b0000000000000001;
        15'b000001111001001 : reciprocal = 16'b0000000000000001;
        15'b000001111001010 : reciprocal = 16'b0000000000000001;
        15'b000001111001011 : reciprocal = 16'b0000000000000001;
        15'b000001111001100 : reciprocal = 16'b0000000000000001;
        15'b000001111001101 : reciprocal = 16'b0000000000000001;
        15'b000001111001110 : reciprocal = 16'b0000000000000001;
        15'b000001111001111 : reciprocal = 16'b0000000000000001;
        15'b000001111010000 : reciprocal = 16'b0000000000000001;
        15'b000001111010001 : reciprocal = 16'b0000000000000001;
        15'b000001111010010 : reciprocal = 16'b0000000000000001;
        15'b000001111010011 : reciprocal = 16'b0000000000000001;
        15'b000001111010100 : reciprocal = 16'b0000000000000001;
        15'b000001111010101 : reciprocal = 16'b0000000000000001;
        15'b000001111010110 : reciprocal = 16'b0000000000000001;
        15'b000001111010111 : reciprocal = 16'b0000000000000001;
        15'b000001111011000 : reciprocal = 16'b0000000000000001;
        15'b000001111011001 : reciprocal = 16'b0000000000000001;
        15'b000001111011010 : reciprocal = 16'b0000000000000001;
        15'b000001111011011 : reciprocal = 16'b0000000000000001;
        15'b000001111011100 : reciprocal = 16'b0000000000000001;
        15'b000001111011101 : reciprocal = 16'b0000000000000001;
        15'b000001111011110 : reciprocal = 16'b0000000000000001;
        15'b000001111011111 : reciprocal = 16'b0000000000000001;
        15'b000001111100000 : reciprocal = 16'b0000000000000001;
        15'b000001111100001 : reciprocal = 16'b0000000000000001;
        15'b000001111100010 : reciprocal = 16'b0000000000000001;
        15'b000001111100011 : reciprocal = 16'b0000000000000001;
        15'b000001111100100 : reciprocal = 16'b0000000000000001;
        15'b000001111100101 : reciprocal = 16'b0000000000000001;
        15'b000001111100110 : reciprocal = 16'b0000000000000001;
        15'b000001111100111 : reciprocal = 16'b0000000000000001;
        15'b000001111101000 : reciprocal = 16'b0000000000000001;
        15'b000001111101001 : reciprocal = 16'b0000000000000001;
        15'b000001111101010 : reciprocal = 16'b0000000000000001;
        15'b000001111101011 : reciprocal = 16'b0000000000000001;
        15'b000001111101100 : reciprocal = 16'b0000000000000001;
        15'b000001111101101 : reciprocal = 16'b0000000000000001;
        15'b000001111101110 : reciprocal = 16'b0000000000000001;
        15'b000001111101111 : reciprocal = 16'b0000000000000001;
        15'b000001111110000 : reciprocal = 16'b0000000000000001;
        15'b000001111110001 : reciprocal = 16'b0000000000000001;
        15'b000001111110010 : reciprocal = 16'b0000000000000001;
        15'b000001111110011 : reciprocal = 16'b0000000000000001;
        15'b000001111110100 : reciprocal = 16'b0000000000000001;
        15'b000001111110101 : reciprocal = 16'b0000000000000001;
        15'b000001111110110 : reciprocal = 16'b0000000000000001;
        15'b000001111110111 : reciprocal = 16'b0000000000000001;
        15'b000001111111000 : reciprocal = 16'b0000000000000001;
        15'b000001111111001 : reciprocal = 16'b0000000000000001;
        15'b000001111111010 : reciprocal = 16'b0000000000000001;
        15'b000001111111011 : reciprocal = 16'b0000000000000001;
        15'b000001111111100 : reciprocal = 16'b0000000000000001;
        15'b000001111111101 : reciprocal = 16'b0000000000000001;
        15'b000001111111110 : reciprocal = 16'b0000000000000001;
        15'b000001111111111 : reciprocal = 16'b0000000000000001;
        default : reciprocal = 16'b0000000000000000;
        15'b111111111111111 : reciprocal = 1111111000000000;
        15'b111111111111110 : reciprocal = 1111111100000000;
        15'b111111111111101 : reciprocal = 1111111101010101;
        15'b111111111111100 : reciprocal = 1111111110000000;
        15'b111111111111011 : reciprocal = 1111111110011010;
        15'b111111111111010 : reciprocal = 1111111110101011;
        15'b111111111111001 : reciprocal = 1111111110110111;
        15'b111111111111000 : reciprocal = 1111111111000000;
        15'b111111111110111 : reciprocal = 1111111111000111;
        15'b111111111110110 : reciprocal = 1111111111001101;
        15'b111111111110101 : reciprocal = 1111111111010001;
        15'b111111111110100 : reciprocal = 1111111111010101;
        15'b111111111110011 : reciprocal = 1111111111011001;
        15'b111111111110010 : reciprocal = 1111111111011011;
        15'b111111111110001 : reciprocal = 1111111111011110;
        15'b111111111110000 : reciprocal = 1111111111100000;
        15'b111111111101111 : reciprocal = 1111111111100010;
        15'b111111111101110 : reciprocal = 1111111111100100;
        15'b111111111101101 : reciprocal = 1111111111100101;
        15'b111111111101100 : reciprocal = 1111111111100110;
        15'b111111111101011 : reciprocal = 1111111111101000;
        15'b111111111101010 : reciprocal = 1111111111101001;
        15'b111111111101001 : reciprocal = 1111111111101010;
        15'b111111111101000 : reciprocal = 1111111111101011;
        15'b111111111100111 : reciprocal = 1111111111101100;
        15'b111111111100110 : reciprocal = 1111111111101100;
        15'b111111111100101 : reciprocal = 1111111111101101;
        15'b111111111100100 : reciprocal = 1111111111101110;
        15'b111111111100011 : reciprocal = 1111111111101110;
        15'b111111111100010 : reciprocal = 1111111111101111;
        15'b111111111100001 : reciprocal = 1111111111101111;
        15'b111111111100000 : reciprocal = 1111111111110000;
        15'b111111111011111 : reciprocal = 1111111111110000;
        15'b111111111011110 : reciprocal = 1111111111110001;
        15'b111111111011101 : reciprocal = 1111111111110001;
        15'b111111111011100 : reciprocal = 1111111111110010;
        15'b111111111011011 : reciprocal = 1111111111110010;
        15'b111111111011010 : reciprocal = 1111111111110011;
        15'b111111111011001 : reciprocal = 1111111111110011;
        15'b111111111011000 : reciprocal = 1111111111110011;
        15'b111111111010111 : reciprocal = 1111111111110100;
        15'b111111111010110 : reciprocal = 1111111111110100;
        15'b111111111010101 : reciprocal = 1111111111110100;
        15'b111111111010100 : reciprocal = 1111111111110100;
        15'b111111111010011 : reciprocal = 1111111111110101;
        15'b111111111010010 : reciprocal = 1111111111110101;
        15'b111111111010001 : reciprocal = 1111111111110101;
        15'b111111111010000 : reciprocal = 1111111111110101;
        15'b111111111001111 : reciprocal = 1111111111110110;
        15'b111111111001110 : reciprocal = 1111111111110110;
        15'b111111111001101 : reciprocal = 1111111111110110;
        15'b111111111001100 : reciprocal = 1111111111110110;
        15'b111111111001011 : reciprocal = 1111111111110110;
        15'b111111111001010 : reciprocal = 1111111111110111;
        15'b111111111001001 : reciprocal = 1111111111110111;
        15'b111111111001000 : reciprocal = 1111111111110111;
        15'b111111111000111 : reciprocal = 1111111111110111;
        15'b111111111000110 : reciprocal = 1111111111110111;
        15'b111111111000101 : reciprocal = 1111111111110111;
        15'b111111111000100 : reciprocal = 1111111111110111;
        15'b111111111000011 : reciprocal = 1111111111111000;
        15'b111111111000010 : reciprocal = 1111111111111000;
        15'b111111111000001 : reciprocal = 1111111111111000;
        15'b111111111000000 : reciprocal = 1111111111111000;
        15'b111111110111111 : reciprocal = 1111111111111000;
        15'b111111110111110 : reciprocal = 1111111111111000;
        15'b111111110111101 : reciprocal = 1111111111111000;
        15'b111111110111100 : reciprocal = 1111111111111000;
        15'b111111110111011 : reciprocal = 1111111111111001;
        15'b111111110111010 : reciprocal = 1111111111111001;
        15'b111111110111001 : reciprocal = 1111111111111001;
        15'b111111110111000 : reciprocal = 1111111111111001;
        15'b111111110110111 : reciprocal = 1111111111111001;
        15'b111111110110110 : reciprocal = 1111111111111001;
        15'b111111110110101 : reciprocal = 1111111111111001;
        15'b111111110110100 : reciprocal = 1111111111111001;
        15'b111111110110011 : reciprocal = 1111111111111001;
        15'b111111110110010 : reciprocal = 1111111111111001;
        15'b111111110110001 : reciprocal = 1111111111111010;
        15'b111111110110000 : reciprocal = 1111111111111010;
        15'b111111110101111 : reciprocal = 1111111111111010;
        15'b111111110101110 : reciprocal = 1111111111111010;
        15'b111111110101101 : reciprocal = 1111111111111010;
        15'b111111110101100 : reciprocal = 1111111111111010;
        15'b111111110101011 : reciprocal = 1111111111111010;
        15'b111111110101010 : reciprocal = 1111111111111010;
        15'b111111110101001 : reciprocal = 1111111111111010;
        15'b111111110101000 : reciprocal = 1111111111111010;
        15'b111111110100111 : reciprocal = 1111111111111010;
        15'b111111110100110 : reciprocal = 1111111111111010;
        15'b111111110100101 : reciprocal = 1111111111111010;
        15'b111111110100100 : reciprocal = 1111111111111010;
        15'b111111110100011 : reciprocal = 1111111111111010;
        15'b111111110100010 : reciprocal = 1111111111111011;
        15'b111111110100001 : reciprocal = 1111111111111011;
        15'b111111110100000 : reciprocal = 1111111111111011;
        15'b111111110011111 : reciprocal = 1111111111111011;
        15'b111111110011110 : reciprocal = 1111111111111011;
        15'b111111110011101 : reciprocal = 1111111111111011;
        15'b111111110011100 : reciprocal = 1111111111111011;
        15'b111111110011011 : reciprocal = 1111111111111011;
        15'b111111110011010 : reciprocal = 1111111111111011;
        15'b111111110011001 : reciprocal = 1111111111111011;
        15'b111111110011000 : reciprocal = 1111111111111011;
        15'b111111110010111 : reciprocal = 1111111111111011;
        15'b111111110010110 : reciprocal = 1111111111111011;
        15'b111111110010101 : reciprocal = 1111111111111011;
        15'b111111110010100 : reciprocal = 1111111111111011;
        15'b111111110010011 : reciprocal = 1111111111111011;
        15'b111111110010010 : reciprocal = 1111111111111011;
        15'b111111110010001 : reciprocal = 1111111111111011;
        15'b111111110010000 : reciprocal = 1111111111111011;
        15'b111111110001111 : reciprocal = 1111111111111011;
        15'b111111110001110 : reciprocal = 1111111111111100;
        15'b111111110001101 : reciprocal = 1111111111111100;
        15'b111111110001100 : reciprocal = 1111111111111100;
        15'b111111110001011 : reciprocal = 1111111111111100;
        15'b111111110001010 : reciprocal = 1111111111111100;
        15'b111111110001001 : reciprocal = 1111111111111100;
        15'b111111110001000 : reciprocal = 1111111111111100;
        15'b111111110000111 : reciprocal = 1111111111111100;
        15'b111111110000110 : reciprocal = 1111111111111100;
        15'b111111110000101 : reciprocal = 1111111111111100;
        15'b111111110000100 : reciprocal = 1111111111111100;
        15'b111111110000011 : reciprocal = 1111111111111100;
        15'b111111110000010 : reciprocal = 1111111111111100;
        15'b111111110000001 : reciprocal = 1111111111111100;
        15'b111111110000000 : reciprocal = 1111111111111100;
        15'b111111101111111 : reciprocal = 1111111111111100;
        15'b111111101111110 : reciprocal = 1111111111111100;
        15'b111111101111101 : reciprocal = 1111111111111100;
        15'b111111101111100 : reciprocal = 1111111111111100;
        15'b111111101111011 : reciprocal = 1111111111111100;
        15'b111111101111010 : reciprocal = 1111111111111100;
        15'b111111101111001 : reciprocal = 1111111111111100;
        15'b111111101111000 : reciprocal = 1111111111111100;
        15'b111111101110111 : reciprocal = 1111111111111100;
        15'b111111101110110 : reciprocal = 1111111111111100;
        15'b111111101110101 : reciprocal = 1111111111111100;
        15'b111111101110100 : reciprocal = 1111111111111100;
        15'b111111101110011 : reciprocal = 1111111111111100;
        15'b111111101110010 : reciprocal = 1111111111111100;
        15'b111111101110001 : reciprocal = 1111111111111100;
        15'b111111101110000 : reciprocal = 1111111111111100;
        15'b111111101101111 : reciprocal = 1111111111111100;
        15'b111111101101110 : reciprocal = 1111111111111100;
        15'b111111101101101 : reciprocal = 1111111111111101;
        15'b111111101101100 : reciprocal = 1111111111111101;
        15'b111111101101011 : reciprocal = 1111111111111101;
        15'b111111101101010 : reciprocal = 1111111111111101;
        15'b111111101101001 : reciprocal = 1111111111111101;
        15'b111111101101000 : reciprocal = 1111111111111101;
        15'b111111101100111 : reciprocal = 1111111111111101;
        15'b111111101100110 : reciprocal = 1111111111111101;
        15'b111111101100101 : reciprocal = 1111111111111101;
        15'b111111101100100 : reciprocal = 1111111111111101;
        15'b111111101100011 : reciprocal = 1111111111111101;
        15'b111111101100010 : reciprocal = 1111111111111101;
        15'b111111101100001 : reciprocal = 1111111111111101;
        15'b111111101100000 : reciprocal = 1111111111111101;
        15'b111111101011111 : reciprocal = 1111111111111101;
        15'b111111101011110 : reciprocal = 1111111111111101;
        15'b111111101011101 : reciprocal = 1111111111111101;
        15'b111111101011100 : reciprocal = 1111111111111101;
        15'b111111101011011 : reciprocal = 1111111111111101;
        15'b111111101011010 : reciprocal = 1111111111111101;
        15'b111111101011001 : reciprocal = 1111111111111101;
        15'b111111101011000 : reciprocal = 1111111111111101;
        15'b111111101010111 : reciprocal = 1111111111111101;
        15'b111111101010110 : reciprocal = 1111111111111101;
        15'b111111101010101 : reciprocal = 1111111111111101;
        15'b111111101010100 : reciprocal = 1111111111111101;
        15'b111111101010011 : reciprocal = 1111111111111101;
        15'b111111101010010 : reciprocal = 1111111111111101;
        15'b111111101010001 : reciprocal = 1111111111111101;
        15'b111111101010000 : reciprocal = 1111111111111101;
        15'b111111101001111 : reciprocal = 1111111111111101;
        15'b111111101001110 : reciprocal = 1111111111111101;
        15'b111111101001101 : reciprocal = 1111111111111101;
        15'b111111101001100 : reciprocal = 1111111111111101;
        15'b111111101001011 : reciprocal = 1111111111111101;
        15'b111111101001010 : reciprocal = 1111111111111101;
        15'b111111101001001 : reciprocal = 1111111111111101;
        15'b111111101001000 : reciprocal = 1111111111111101;
        15'b111111101000111 : reciprocal = 1111111111111101;
        15'b111111101000110 : reciprocal = 1111111111111101;
        15'b111111101000101 : reciprocal = 1111111111111101;
        15'b111111101000100 : reciprocal = 1111111111111101;
        15'b111111101000011 : reciprocal = 1111111111111101;
        15'b111111101000010 : reciprocal = 1111111111111101;
        15'b111111101000001 : reciprocal = 1111111111111101;
        15'b111111101000000 : reciprocal = 1111111111111101;
        15'b111111100111111 : reciprocal = 1111111111111101;
        15'b111111100111110 : reciprocal = 1111111111111101;
        15'b111111100111101 : reciprocal = 1111111111111101;
        15'b111111100111100 : reciprocal = 1111111111111101;
        15'b111111100111011 : reciprocal = 1111111111111101;
        15'b111111100111010 : reciprocal = 1111111111111101;
        15'b111111100111001 : reciprocal = 1111111111111101;
        15'b111111100111000 : reciprocal = 1111111111111101;
        15'b111111100110111 : reciprocal = 1111111111111101;
        15'b111111100110110 : reciprocal = 1111111111111101;
        15'b111111100110101 : reciprocal = 1111111111111101;
        15'b111111100110100 : reciprocal = 1111111111111101;
        15'b111111100110011 : reciprocal = 1111111111111110;
        15'b111111100110010 : reciprocal = 1111111111111110;
        15'b111111100110001 : reciprocal = 1111111111111110;
        15'b111111100110000 : reciprocal = 1111111111111110;
        15'b111111100101111 : reciprocal = 1111111111111110;
        15'b111111100101110 : reciprocal = 1111111111111110;
        15'b111111100101101 : reciprocal = 1111111111111110;
        15'b111111100101100 : reciprocal = 1111111111111110;
        15'b111111100101011 : reciprocal = 1111111111111110;
        15'b111111100101010 : reciprocal = 1111111111111110;
        15'b111111100101001 : reciprocal = 1111111111111110;
        15'b111111100101000 : reciprocal = 1111111111111110;
        15'b111111100100111 : reciprocal = 1111111111111110;
        15'b111111100100110 : reciprocal = 1111111111111110;
        15'b111111100100101 : reciprocal = 1111111111111110;
        15'b111111100100100 : reciprocal = 1111111111111110;
        15'b111111100100011 : reciprocal = 1111111111111110;
        15'b111111100100010 : reciprocal = 1111111111111110;
        15'b111111100100001 : reciprocal = 1111111111111110;
        15'b111111100100000 : reciprocal = 1111111111111110;
        15'b111111100011111 : reciprocal = 1111111111111110;
        15'b111111100011110 : reciprocal = 1111111111111110;
        15'b111111100011101 : reciprocal = 1111111111111110;
        15'b111111100011100 : reciprocal = 1111111111111110;
        15'b111111100011011 : reciprocal = 1111111111111110;
        15'b111111100011010 : reciprocal = 1111111111111110;
        15'b111111100011001 : reciprocal = 1111111111111110;
        15'b111111100011000 : reciprocal = 1111111111111110;
        15'b111111100010111 : reciprocal = 1111111111111110;
        15'b111111100010110 : reciprocal = 1111111111111110;
        15'b111111100010101 : reciprocal = 1111111111111110;
        15'b111111100010100 : reciprocal = 1111111111111110;
        15'b111111100010011 : reciprocal = 1111111111111110;
        15'b111111100010010 : reciprocal = 1111111111111110;
        15'b111111100010001 : reciprocal = 1111111111111110;
        15'b111111100010000 : reciprocal = 1111111111111110;
        15'b111111100001111 : reciprocal = 1111111111111110;
        15'b111111100001110 : reciprocal = 1111111111111110;
        15'b111111100001101 : reciprocal = 1111111111111110;
        15'b111111100001100 : reciprocal = 1111111111111110;
        15'b111111100001011 : reciprocal = 1111111111111110;
        15'b111111100001010 : reciprocal = 1111111111111110;
        15'b111111100001001 : reciprocal = 1111111111111110;
        15'b111111100001000 : reciprocal = 1111111111111110;
        15'b111111100000111 : reciprocal = 1111111111111110;
        15'b111111100000110 : reciprocal = 1111111111111110;
        15'b111111100000101 : reciprocal = 1111111111111110;
        15'b111111100000100 : reciprocal = 1111111111111110;
        15'b111111100000011 : reciprocal = 1111111111111110;
        15'b111111100000010 : reciprocal = 1111111111111110;
        15'b111111100000001 : reciprocal = 1111111111111110;
        15'b111111100000000 : reciprocal = 1111111111111110;
        15'b111111011111111 : reciprocal = 1111111111111110;
        15'b111111011111110 : reciprocal = 1111111111111110;
        15'b111111011111101 : reciprocal = 1111111111111110;
        15'b111111011111100 : reciprocal = 1111111111111110;
        15'b111111011111011 : reciprocal = 1111111111111110;
        15'b111111011111010 : reciprocal = 1111111111111110;
        15'b111111011111001 : reciprocal = 1111111111111110;
        15'b111111011111000 : reciprocal = 1111111111111110;
        15'b111111011110111 : reciprocal = 1111111111111110;
        15'b111111011110110 : reciprocal = 1111111111111110;
        15'b111111011110101 : reciprocal = 1111111111111110;
        15'b111111011110100 : reciprocal = 1111111111111110;
        15'b111111011110011 : reciprocal = 1111111111111110;
        15'b111111011110010 : reciprocal = 1111111111111110;
        15'b111111011110001 : reciprocal = 1111111111111110;
        15'b111111011110000 : reciprocal = 1111111111111110;
        15'b111111011101111 : reciprocal = 1111111111111110;
        15'b111111011101110 : reciprocal = 1111111111111110;
        15'b111111011101101 : reciprocal = 1111111111111110;
        15'b111111011101100 : reciprocal = 1111111111111110;
        15'b111111011101011 : reciprocal = 1111111111111110;
        15'b111111011101010 : reciprocal = 1111111111111110;
        15'b111111011101001 : reciprocal = 1111111111111110;
        15'b111111011101000 : reciprocal = 1111111111111110;
        15'b111111011100111 : reciprocal = 1111111111111110;
        15'b111111011100110 : reciprocal = 1111111111111110;
        15'b111111011100101 : reciprocal = 1111111111111110;
        15'b111111011100100 : reciprocal = 1111111111111110;
        15'b111111011100011 : reciprocal = 1111111111111110;
        15'b111111011100010 : reciprocal = 1111111111111110;
        15'b111111011100001 : reciprocal = 1111111111111110;
        15'b111111011100000 : reciprocal = 1111111111111110;
        15'b111111011011111 : reciprocal = 1111111111111110;
        15'b111111011011110 : reciprocal = 1111111111111110;
        15'b111111011011101 : reciprocal = 1111111111111110;
        15'b111111011011100 : reciprocal = 1111111111111110;
        15'b111111011011011 : reciprocal = 1111111111111110;
        15'b111111011011010 : reciprocal = 1111111111111110;
        15'b111111011011001 : reciprocal = 1111111111111110;
        15'b111111011011000 : reciprocal = 1111111111111110;
        15'b111111011010111 : reciprocal = 1111111111111110;
        15'b111111011010110 : reciprocal = 1111111111111110;
        15'b111111011010101 : reciprocal = 1111111111111110;
        15'b111111011010100 : reciprocal = 1111111111111110;
        15'b111111011010011 : reciprocal = 1111111111111110;
        15'b111111011010010 : reciprocal = 1111111111111110;
        15'b111111011010001 : reciprocal = 1111111111111110;
        15'b111111011010000 : reciprocal = 1111111111111110;
        15'b111111011001111 : reciprocal = 1111111111111110;
        15'b111111011001110 : reciprocal = 1111111111111110;
        15'b111111011001101 : reciprocal = 1111111111111110;
        15'b111111011001100 : reciprocal = 1111111111111110;
        15'b111111011001011 : reciprocal = 1111111111111110;
        15'b111111011001010 : reciprocal = 1111111111111110;
        15'b111111011001001 : reciprocal = 1111111111111110;
        15'b111111011001000 : reciprocal = 1111111111111110;
        15'b111111011000111 : reciprocal = 1111111111111110;
        15'b111111011000110 : reciprocal = 1111111111111110;
        15'b111111011000101 : reciprocal = 1111111111111110;
        15'b111111011000100 : reciprocal = 1111111111111110;
        15'b111111011000011 : reciprocal = 1111111111111110;
        15'b111111011000010 : reciprocal = 1111111111111110;
        15'b111111011000001 : reciprocal = 1111111111111110;
        15'b111111011000000 : reciprocal = 1111111111111110;
        15'b111111010111111 : reciprocal = 1111111111111110;
        15'b111111010111110 : reciprocal = 1111111111111110;
        15'b111111010111101 : reciprocal = 1111111111111110;
        15'b111111010111100 : reciprocal = 1111111111111110;
        15'b111111010111011 : reciprocal = 1111111111111110;
        15'b111111010111010 : reciprocal = 1111111111111110;
        15'b111111010111001 : reciprocal = 1111111111111110;
        15'b111111010111000 : reciprocal = 1111111111111110;
        15'b111111010110111 : reciprocal = 1111111111111110;
        15'b111111010110110 : reciprocal = 1111111111111110;
        15'b111111010110101 : reciprocal = 1111111111111110;
        15'b111111010110100 : reciprocal = 1111111111111110;
        15'b111111010110011 : reciprocal = 1111111111111110;
        15'b111111010110010 : reciprocal = 1111111111111110;
        15'b111111010110001 : reciprocal = 1111111111111110;
        15'b111111010110000 : reciprocal = 1111111111111110;
        15'b111111010101111 : reciprocal = 1111111111111110;
        15'b111111010101110 : reciprocal = 1111111111111110;
        15'b111111010101101 : reciprocal = 1111111111111110;
        15'b111111010101100 : reciprocal = 1111111111111110;
        15'b111111010101011 : reciprocal = 1111111111111110;
        15'b111111010101010 : reciprocal = 1111111111111111;
        15'b111111010101001 : reciprocal = 1111111111111111;
        15'b111111010101000 : reciprocal = 1111111111111111;
        15'b111111010100111 : reciprocal = 1111111111111111;
        15'b111111010100110 : reciprocal = 1111111111111111;
        15'b111111010100101 : reciprocal = 1111111111111111;
        15'b111111010100100 : reciprocal = 1111111111111111;
        15'b111111010100011 : reciprocal = 1111111111111111;
        15'b111111010100010 : reciprocal = 1111111111111111;
        15'b111111010100001 : reciprocal = 1111111111111111;
        15'b111111010100000 : reciprocal = 1111111111111111;
        15'b111111010011111 : reciprocal = 1111111111111111;
        15'b111111010011110 : reciprocal = 1111111111111111;
        15'b111111010011101 : reciprocal = 1111111111111111;
        15'b111111010011100 : reciprocal = 1111111111111111;
        15'b111111010011011 : reciprocal = 1111111111111111;
        15'b111111010011010 : reciprocal = 1111111111111111;
        15'b111111010011001 : reciprocal = 1111111111111111;
        15'b111111010011000 : reciprocal = 1111111111111111;
        15'b111111010010111 : reciprocal = 1111111111111111;
        15'b111111010010110 : reciprocal = 1111111111111111;
        15'b111111010010101 : reciprocal = 1111111111111111;
        15'b111111010010100 : reciprocal = 1111111111111111;
        15'b111111010010011 : reciprocal = 1111111111111111;
        15'b111111010010010 : reciprocal = 1111111111111111;
        15'b111111010010001 : reciprocal = 1111111111111111;
        15'b111111010010000 : reciprocal = 1111111111111111;
        15'b111111010001111 : reciprocal = 1111111111111111;
        15'b111111010001110 : reciprocal = 1111111111111111;
        15'b111111010001101 : reciprocal = 1111111111111111;
        15'b111111010001100 : reciprocal = 1111111111111111;
        15'b111111010001011 : reciprocal = 1111111111111111;
        15'b111111010001010 : reciprocal = 1111111111111111;
        15'b111111010001001 : reciprocal = 1111111111111111;
        15'b111111010001000 : reciprocal = 1111111111111111;
        15'b111111010000111 : reciprocal = 1111111111111111;
        15'b111111010000110 : reciprocal = 1111111111111111;
        15'b111111010000101 : reciprocal = 1111111111111111;
        15'b111111010000100 : reciprocal = 1111111111111111;
        15'b111111010000011 : reciprocal = 1111111111111111;
        15'b111111010000010 : reciprocal = 1111111111111111;
        15'b111111010000001 : reciprocal = 1111111111111111;
        15'b111111010000000 : reciprocal = 1111111111111111;
        15'b111111001111111 : reciprocal = 1111111111111111;
        15'b111111001111110 : reciprocal = 1111111111111111;
        15'b111111001111101 : reciprocal = 1111111111111111;
        15'b111111001111100 : reciprocal = 1111111111111111;
        15'b111111001111011 : reciprocal = 1111111111111111;
        15'b111111001111010 : reciprocal = 1111111111111111;
        15'b111111001111001 : reciprocal = 1111111111111111;
        15'b111111001111000 : reciprocal = 1111111111111111;
        15'b111111001110111 : reciprocal = 1111111111111111;
        15'b111111001110110 : reciprocal = 1111111111111111;
        15'b111111001110101 : reciprocal = 1111111111111111;
        15'b111111001110100 : reciprocal = 1111111111111111;
        15'b111111001110011 : reciprocal = 1111111111111111;
        15'b111111001110010 : reciprocal = 1111111111111111;
        15'b111111001110001 : reciprocal = 1111111111111111;
        15'b111111001110000 : reciprocal = 1111111111111111;
        15'b111111001101111 : reciprocal = 1111111111111111;
        15'b111111001101110 : reciprocal = 1111111111111111;
        15'b111111001101101 : reciprocal = 1111111111111111;
        15'b111111001101100 : reciprocal = 1111111111111111;
        15'b111111001101011 : reciprocal = 1111111111111111;
        15'b111111001101010 : reciprocal = 1111111111111111;
        15'b111111001101001 : reciprocal = 1111111111111111;
        15'b111111001101000 : reciprocal = 1111111111111111;
        15'b111111001100111 : reciprocal = 1111111111111111;
        15'b111111001100110 : reciprocal = 1111111111111111;
        15'b111111001100101 : reciprocal = 1111111111111111;
        15'b111111001100100 : reciprocal = 1111111111111111;
        15'b111111001100011 : reciprocal = 1111111111111111;
        15'b111111001100010 : reciprocal = 1111111111111111;
        15'b111111001100001 : reciprocal = 1111111111111111;
        15'b111111001100000 : reciprocal = 1111111111111111;
        15'b111111001011111 : reciprocal = 1111111111111111;
        15'b111111001011110 : reciprocal = 1111111111111111;
        15'b111111001011101 : reciprocal = 1111111111111111;
        15'b111111001011100 : reciprocal = 1111111111111111;
        15'b111111001011011 : reciprocal = 1111111111111111;
        15'b111111001011010 : reciprocal = 1111111111111111;
        15'b111111001011001 : reciprocal = 1111111111111111;
        15'b111111001011000 : reciprocal = 1111111111111111;
        15'b111111001010111 : reciprocal = 1111111111111111;
        15'b111111001010110 : reciprocal = 1111111111111111;
        15'b111111001010101 : reciprocal = 1111111111111111;
        15'b111111001010100 : reciprocal = 1111111111111111;
        15'b111111001010011 : reciprocal = 1111111111111111;
        15'b111111001010010 : reciprocal = 1111111111111111;
        15'b111111001010001 : reciprocal = 1111111111111111;
        15'b111111001010000 : reciprocal = 1111111111111111;
        15'b111111001001111 : reciprocal = 1111111111111111;
        15'b111111001001110 : reciprocal = 1111111111111111;
        15'b111111001001101 : reciprocal = 1111111111111111;
        15'b111111001001100 : reciprocal = 1111111111111111;
        15'b111111001001011 : reciprocal = 1111111111111111;
        15'b111111001001010 : reciprocal = 1111111111111111;
        15'b111111001001001 : reciprocal = 1111111111111111;
        15'b111111001001000 : reciprocal = 1111111111111111;
        15'b111111001000111 : reciprocal = 1111111111111111;
        15'b111111001000110 : reciprocal = 1111111111111111;
        15'b111111001000101 : reciprocal = 1111111111111111;
        15'b111111001000100 : reciprocal = 1111111111111111;
        15'b111111001000011 : reciprocal = 1111111111111111;
        15'b111111001000010 : reciprocal = 1111111111111111;
        15'b111111001000001 : reciprocal = 1111111111111111;
        15'b111111001000000 : reciprocal = 1111111111111111;
        15'b111111000111111 : reciprocal = 1111111111111111;
        15'b111111000111110 : reciprocal = 1111111111111111;
        15'b111111000111101 : reciprocal = 1111111111111111;
        15'b111111000111100 : reciprocal = 1111111111111111;
        15'b111111000111011 : reciprocal = 1111111111111111;
        15'b111111000111010 : reciprocal = 1111111111111111;
        15'b111111000111001 : reciprocal = 1111111111111111;
        15'b111111000111000 : reciprocal = 1111111111111111;
        15'b111111000110111 : reciprocal = 1111111111111111;
        15'b111111000110110 : reciprocal = 1111111111111111;
        15'b111111000110101 : reciprocal = 1111111111111111;
        15'b111111000110100 : reciprocal = 1111111111111111;
        15'b111111000110011 : reciprocal = 1111111111111111;
        15'b111111000110010 : reciprocal = 1111111111111111;
        15'b111111000110001 : reciprocal = 1111111111111111;
        15'b111111000110000 : reciprocal = 1111111111111111;
        15'b111111000101111 : reciprocal = 1111111111111111;
        15'b111111000101110 : reciprocal = 1111111111111111;
        15'b111111000101101 : reciprocal = 1111111111111111;
        15'b111111000101100 : reciprocal = 1111111111111111;
        15'b111111000101011 : reciprocal = 1111111111111111;
        15'b111111000101010 : reciprocal = 1111111111111111;
        15'b111111000101001 : reciprocal = 1111111111111111;
        15'b111111000101000 : reciprocal = 1111111111111111;
        15'b111111000100111 : reciprocal = 1111111111111111;
        15'b111111000100110 : reciprocal = 1111111111111111;
        15'b111111000100101 : reciprocal = 1111111111111111;
        15'b111111000100100 : reciprocal = 1111111111111111;
        15'b111111000100011 : reciprocal = 1111111111111111;
        15'b111111000100010 : reciprocal = 1111111111111111;
        15'b111111000100001 : reciprocal = 1111111111111111;
        15'b111111000100000 : reciprocal = 1111111111111111;
        15'b111111000011111 : reciprocal = 1111111111111111;
        15'b111111000011110 : reciprocal = 1111111111111111;
        15'b111111000011101 : reciprocal = 1111111111111111;
        15'b111111000011100 : reciprocal = 1111111111111111;
        15'b111111000011011 : reciprocal = 1111111111111111;
        15'b111111000011010 : reciprocal = 1111111111111111;
        15'b111111000011001 : reciprocal = 1111111111111111;
        15'b111111000011000 : reciprocal = 1111111111111111;
        15'b111111000010111 : reciprocal = 1111111111111111;
        15'b111111000010110 : reciprocal = 1111111111111111;
        15'b111111000010101 : reciprocal = 1111111111111111;
        15'b111111000010100 : reciprocal = 1111111111111111;
        15'b111111000010011 : reciprocal = 1111111111111111;
        15'b111111000010010 : reciprocal = 1111111111111111;
        15'b111111000010001 : reciprocal = 1111111111111111;
        15'b111111000010000 : reciprocal = 1111111111111111;
        15'b111111000001111 : reciprocal = 1111111111111111;
        15'b111111000001110 : reciprocal = 1111111111111111;
        15'b111111000001101 : reciprocal = 1111111111111111;
        15'b111111000001100 : reciprocal = 1111111111111111;
        15'b111111000001011 : reciprocal = 1111111111111111;
        15'b111111000001010 : reciprocal = 1111111111111111;
        15'b111111000001001 : reciprocal = 1111111111111111;
        15'b111111000001000 : reciprocal = 1111111111111111;
        15'b111111000000111 : reciprocal = 1111111111111111;
        15'b111111000000110 : reciprocal = 1111111111111111;
        15'b111111000000101 : reciprocal = 1111111111111111;
        15'b111111000000100 : reciprocal = 1111111111111111;
        15'b111111000000011 : reciprocal = 1111111111111111;
        15'b111111000000010 : reciprocal = 1111111111111111;
        15'b111111000000001 : reciprocal = 1111111111111111;
        15'b111111000000000 : reciprocal = 1111111111111111;
        15'b111110111111111 : reciprocal = 1111111111111111;
        15'b111110111111110 : reciprocal = 1111111111111111;
        15'b111110111111101 : reciprocal = 1111111111111111;
        15'b111110111111100 : reciprocal = 1111111111111111;
        15'b111110111111011 : reciprocal = 1111111111111111;
        15'b111110111111010 : reciprocal = 1111111111111111;
        15'b111110111111001 : reciprocal = 1111111111111111;
        15'b111110111111000 : reciprocal = 1111111111111111;
        15'b111110111110111 : reciprocal = 1111111111111111;
        15'b111110111110110 : reciprocal = 1111111111111111;
        15'b111110111110101 : reciprocal = 1111111111111111;
        15'b111110111110100 : reciprocal = 1111111111111111;
        15'b111110111110011 : reciprocal = 1111111111111111;
        15'b111110111110010 : reciprocal = 1111111111111111;
        15'b111110111110001 : reciprocal = 1111111111111111;
        15'b111110111110000 : reciprocal = 1111111111111111;
        15'b111110111101111 : reciprocal = 1111111111111111;
        15'b111110111101110 : reciprocal = 1111111111111111;
        15'b111110111101101 : reciprocal = 1111111111111111;
        15'b111110111101100 : reciprocal = 1111111111111111;
        15'b111110111101011 : reciprocal = 1111111111111111;
        15'b111110111101010 : reciprocal = 1111111111111111;
        15'b111110111101001 : reciprocal = 1111111111111111;
        15'b111110111101000 : reciprocal = 1111111111111111;
        15'b111110111100111 : reciprocal = 1111111111111111;
        15'b111110111100110 : reciprocal = 1111111111111111;
        15'b111110111100101 : reciprocal = 1111111111111111;
        15'b111110111100100 : reciprocal = 1111111111111111;
        15'b111110111100011 : reciprocal = 1111111111111111;
        15'b111110111100010 : reciprocal = 1111111111111111;
        15'b111110111100001 : reciprocal = 1111111111111111;
        15'b111110111100000 : reciprocal = 1111111111111111;
        15'b111110111011111 : reciprocal = 1111111111111111;
        15'b111110111011110 : reciprocal = 1111111111111111;
        15'b111110111011101 : reciprocal = 1111111111111111;
        15'b111110111011100 : reciprocal = 1111111111111111;
        15'b111110111011011 : reciprocal = 1111111111111111;
        15'b111110111011010 : reciprocal = 1111111111111111;
        15'b111110111011001 : reciprocal = 1111111111111111;
        15'b111110111011000 : reciprocal = 1111111111111111;
        15'b111110111010111 : reciprocal = 1111111111111111;
        15'b111110111010110 : reciprocal = 1111111111111111;
        15'b111110111010101 : reciprocal = 1111111111111111;
        15'b111110111010100 : reciprocal = 1111111111111111;
        15'b111110111010011 : reciprocal = 1111111111111111;
        15'b111110111010010 : reciprocal = 1111111111111111;
        15'b111110111010001 : reciprocal = 1111111111111111;
        15'b111110111010000 : reciprocal = 1111111111111111;
        15'b111110111001111 : reciprocal = 1111111111111111;
        15'b111110111001110 : reciprocal = 1111111111111111;
        15'b111110111001101 : reciprocal = 1111111111111111;
        15'b111110111001100 : reciprocal = 1111111111111111;
        15'b111110111001011 : reciprocal = 1111111111111111;
        15'b111110111001010 : reciprocal = 1111111111111111;
        15'b111110111001001 : reciprocal = 1111111111111111;
        15'b111110111001000 : reciprocal = 1111111111111111;
        15'b111110111000111 : reciprocal = 1111111111111111;
        15'b111110111000110 : reciprocal = 1111111111111111;
        15'b111110111000101 : reciprocal = 1111111111111111;
        15'b111110111000100 : reciprocal = 1111111111111111;
        15'b111110111000011 : reciprocal = 1111111111111111;
        15'b111110111000010 : reciprocal = 1111111111111111;
        15'b111110111000001 : reciprocal = 1111111111111111;
        15'b111110111000000 : reciprocal = 1111111111111111;
        15'b111110110111111 : reciprocal = 1111111111111111;
        15'b111110110111110 : reciprocal = 1111111111111111;
        15'b111110110111101 : reciprocal = 1111111111111111;
        15'b111110110111100 : reciprocal = 1111111111111111;
        15'b111110110111011 : reciprocal = 1111111111111111;
        15'b111110110111010 : reciprocal = 1111111111111111;
        15'b111110110111001 : reciprocal = 1111111111111111;
        15'b111110110111000 : reciprocal = 1111111111111111;
        15'b111110110110111 : reciprocal = 1111111111111111;
        15'b111110110110110 : reciprocal = 1111111111111111;
        15'b111110110110101 : reciprocal = 1111111111111111;
        15'b111110110110100 : reciprocal = 1111111111111111;
        15'b111110110110011 : reciprocal = 1111111111111111;
        15'b111110110110010 : reciprocal = 1111111111111111;
        15'b111110110110001 : reciprocal = 1111111111111111;
        15'b111110110110000 : reciprocal = 1111111111111111;
        15'b111110110101111 : reciprocal = 1111111111111111;
        15'b111110110101110 : reciprocal = 1111111111111111;
        15'b111110110101101 : reciprocal = 1111111111111111;
        15'b111110110101100 : reciprocal = 1111111111111111;
        15'b111110110101011 : reciprocal = 1111111111111111;
        15'b111110110101010 : reciprocal = 1111111111111111;
        15'b111110110101001 : reciprocal = 1111111111111111;
        15'b111110110101000 : reciprocal = 1111111111111111;
        15'b111110110100111 : reciprocal = 1111111111111111;
        15'b111110110100110 : reciprocal = 1111111111111111;
        15'b111110110100101 : reciprocal = 1111111111111111;
        15'b111110110100100 : reciprocal = 1111111111111111;
        15'b111110110100011 : reciprocal = 1111111111111111;
        15'b111110110100010 : reciprocal = 1111111111111111;
        15'b111110110100001 : reciprocal = 1111111111111111;
        15'b111110110100000 : reciprocal = 1111111111111111;
        15'b111110110011111 : reciprocal = 1111111111111111;
        15'b111110110011110 : reciprocal = 1111111111111111;
        15'b111110110011101 : reciprocal = 1111111111111111;
        15'b111110110011100 : reciprocal = 1111111111111111;
        15'b111110110011011 : reciprocal = 1111111111111111;
        15'b111110110011010 : reciprocal = 1111111111111111;
        15'b111110110011001 : reciprocal = 1111111111111111;
        15'b111110110011000 : reciprocal = 1111111111111111;
        15'b111110110010111 : reciprocal = 1111111111111111;
        15'b111110110010110 : reciprocal = 1111111111111111;
        15'b111110110010101 : reciprocal = 1111111111111111;
        15'b111110110010100 : reciprocal = 1111111111111111;
        15'b111110110010011 : reciprocal = 1111111111111111;
        15'b111110110010010 : reciprocal = 1111111111111111;
        15'b111110110010001 : reciprocal = 1111111111111111;
        15'b111110110010000 : reciprocal = 1111111111111111;
        15'b111110110001111 : reciprocal = 1111111111111111;
        15'b111110110001110 : reciprocal = 1111111111111111;
        15'b111110110001101 : reciprocal = 1111111111111111;
        15'b111110110001100 : reciprocal = 1111111111111111;
        15'b111110110001011 : reciprocal = 1111111111111111;
        15'b111110110001010 : reciprocal = 1111111111111111;
        15'b111110110001001 : reciprocal = 1111111111111111;
        15'b111110110001000 : reciprocal = 1111111111111111;
        15'b111110110000111 : reciprocal = 1111111111111111;
        15'b111110110000110 : reciprocal = 1111111111111111;
        15'b111110110000101 : reciprocal = 1111111111111111;
        15'b111110110000100 : reciprocal = 1111111111111111;
        15'b111110110000011 : reciprocal = 1111111111111111;
        15'b111110110000010 : reciprocal = 1111111111111111;
        15'b111110110000001 : reciprocal = 1111111111111111;
        15'b111110110000000 : reciprocal = 1111111111111111;
        15'b111110101111111 : reciprocal = 1111111111111111;
        15'b111110101111110 : reciprocal = 1111111111111111;
        15'b111110101111101 : reciprocal = 1111111111111111;
        15'b111110101111100 : reciprocal = 1111111111111111;
        15'b111110101111011 : reciprocal = 1111111111111111;
        15'b111110101111010 : reciprocal = 1111111111111111;
        15'b111110101111001 : reciprocal = 1111111111111111;
        15'b111110101111000 : reciprocal = 1111111111111111;
        15'b111110101110111 : reciprocal = 1111111111111111;
        15'b111110101110110 : reciprocal = 1111111111111111;
        15'b111110101110101 : reciprocal = 1111111111111111;
        15'b111110101110100 : reciprocal = 1111111111111111;
        15'b111110101110011 : reciprocal = 1111111111111111;
        15'b111110101110010 : reciprocal = 1111111111111111;
        15'b111110101110001 : reciprocal = 1111111111111111;
        15'b111110101110000 : reciprocal = 1111111111111111;
        15'b111110101101111 : reciprocal = 1111111111111111;
        15'b111110101101110 : reciprocal = 1111111111111111;
        15'b111110101101101 : reciprocal = 1111111111111111;
        15'b111110101101100 : reciprocal = 1111111111111111;
        15'b111110101101011 : reciprocal = 1111111111111111;
        15'b111110101101010 : reciprocal = 1111111111111111;
        15'b111110101101001 : reciprocal = 1111111111111111;
        15'b111110101101000 : reciprocal = 1111111111111111;
        15'b111110101100111 : reciprocal = 1111111111111111;
        15'b111110101100110 : reciprocal = 1111111111111111;
        15'b111110101100101 : reciprocal = 1111111111111111;
        15'b111110101100100 : reciprocal = 1111111111111111;
        15'b111110101100011 : reciprocal = 1111111111111111;
        15'b111110101100010 : reciprocal = 1111111111111111;
        15'b111110101100001 : reciprocal = 1111111111111111;
        15'b111110101100000 : reciprocal = 1111111111111111;
        15'b111110101011111 : reciprocal = 1111111111111111;
        15'b111110101011110 : reciprocal = 1111111111111111;
        15'b111110101011101 : reciprocal = 1111111111111111;
        15'b111110101011100 : reciprocal = 1111111111111111;
        15'b111110101011011 : reciprocal = 1111111111111111;
        15'b111110101011010 : reciprocal = 1111111111111111;
        15'b111110101011001 : reciprocal = 1111111111111111;
        15'b111110101011000 : reciprocal = 1111111111111111;
        15'b111110101010111 : reciprocal = 1111111111111111;
        15'b111110101010110 : reciprocal = 1111111111111111;
        15'b111110101010101 : reciprocal = 1111111111111111;
        15'b111110101010100 : reciprocal = 1111111111111111;
        15'b111110101010011 : reciprocal = 1111111111111111;
        15'b111110101010010 : reciprocal = 1111111111111111;
        15'b111110101010001 : reciprocal = 1111111111111111;
        15'b111110101010000 : reciprocal = 1111111111111111;
        15'b111110101001111 : reciprocal = 1111111111111111;
        15'b111110101001110 : reciprocal = 1111111111111111;
        15'b111110101001101 : reciprocal = 1111111111111111;
        15'b111110101001100 : reciprocal = 1111111111111111;
        15'b111110101001011 : reciprocal = 1111111111111111;
        15'b111110101001010 : reciprocal = 1111111111111111;
        15'b111110101001001 : reciprocal = 1111111111111111;
        15'b111110101001000 : reciprocal = 1111111111111111;
        15'b111110101000111 : reciprocal = 1111111111111111;
        15'b111110101000110 : reciprocal = 1111111111111111;
        15'b111110101000101 : reciprocal = 1111111111111111;
        15'b111110101000100 : reciprocal = 1111111111111111;
        15'b111110101000011 : reciprocal = 1111111111111111;
        15'b111110101000010 : reciprocal = 1111111111111111;
        15'b111110101000001 : reciprocal = 1111111111111111;
        15'b111110101000000 : reciprocal = 1111111111111111;
        15'b111110100111111 : reciprocal = 1111111111111111;
        15'b111110100111110 : reciprocal = 1111111111111111;
        15'b111110100111101 : reciprocal = 1111111111111111;
        15'b111110100111100 : reciprocal = 1111111111111111;
        15'b111110100111011 : reciprocal = 1111111111111111;
        15'b111110100111010 : reciprocal = 1111111111111111;
        15'b111110100111001 : reciprocal = 1111111111111111;
        15'b111110100111000 : reciprocal = 1111111111111111;
        15'b111110100110111 : reciprocal = 1111111111111111;
        15'b111110100110110 : reciprocal = 1111111111111111;
        15'b111110100110101 : reciprocal = 1111111111111111;
        15'b111110100110100 : reciprocal = 1111111111111111;
        15'b111110100110011 : reciprocal = 1111111111111111;
        15'b111110100110010 : reciprocal = 1111111111111111;
        15'b111110100110001 : reciprocal = 1111111111111111;
        15'b111110100110000 : reciprocal = 1111111111111111;
        15'b111110100101111 : reciprocal = 1111111111111111;
        15'b111110100101110 : reciprocal = 1111111111111111;
        15'b111110100101101 : reciprocal = 1111111111111111;
        15'b111110100101100 : reciprocal = 1111111111111111;
        15'b111110100101011 : reciprocal = 1111111111111111;
        15'b111110100101010 : reciprocal = 1111111111111111;
        15'b111110100101001 : reciprocal = 1111111111111111;
        15'b111110100101000 : reciprocal = 1111111111111111;
        15'b111110100100111 : reciprocal = 1111111111111111;
        15'b111110100100110 : reciprocal = 1111111111111111;
        15'b111110100100101 : reciprocal = 1111111111111111;
        15'b111110100100100 : reciprocal = 1111111111111111;
        15'b111110100100011 : reciprocal = 1111111111111111;
        15'b111110100100010 : reciprocal = 1111111111111111;
        15'b111110100100001 : reciprocal = 1111111111111111;
        15'b111110100100000 : reciprocal = 1111111111111111;
        15'b111110100011111 : reciprocal = 1111111111111111;
        15'b111110100011110 : reciprocal = 1111111111111111;
        15'b111110100011101 : reciprocal = 1111111111111111;
        15'b111110100011100 : reciprocal = 1111111111111111;
        15'b111110100011011 : reciprocal = 1111111111111111;
        15'b111110100011010 : reciprocal = 1111111111111111;
        15'b111110100011001 : reciprocal = 1111111111111111;
        15'b111110100011000 : reciprocal = 1111111111111111;
        15'b111110100010111 : reciprocal = 1111111111111111;
        15'b111110100010110 : reciprocal = 1111111111111111;
        15'b111110100010101 : reciprocal = 1111111111111111;
        15'b111110100010100 : reciprocal = 1111111111111111;
        15'b111110100010011 : reciprocal = 1111111111111111;
        15'b111110100010010 : reciprocal = 1111111111111111;
        15'b111110100010001 : reciprocal = 1111111111111111;
        15'b111110100010000 : reciprocal = 1111111111111111;
        15'b111110100001111 : reciprocal = 1111111111111111;
        15'b111110100001110 : reciprocal = 1111111111111111;
        15'b111110100001101 : reciprocal = 1111111111111111;
        15'b111110100001100 : reciprocal = 1111111111111111;
        15'b111110100001011 : reciprocal = 1111111111111111;
        15'b111110100001010 : reciprocal = 1111111111111111;
        15'b111110100001001 : reciprocal = 1111111111111111;
        15'b111110100001000 : reciprocal = 1111111111111111;
        15'b111110100000111 : reciprocal = 1111111111111111;
        15'b111110100000110 : reciprocal = 1111111111111111;
        15'b111110100000101 : reciprocal = 1111111111111111;
        15'b111110100000100 : reciprocal = 1111111111111111;
        15'b111110100000011 : reciprocal = 1111111111111111;
        15'b111110100000010 : reciprocal = 1111111111111111;
        15'b111110100000001 : reciprocal = 1111111111111111;
        15'b111110100000000 : reciprocal = 1111111111111111;
        15'b111110011111111 : reciprocal = 1111111111111111;
        15'b111110011111110 : reciprocal = 1111111111111111;
        15'b111110011111101 : reciprocal = 1111111111111111;
        15'b111110011111100 : reciprocal = 1111111111111111;
        15'b111110011111011 : reciprocal = 1111111111111111;
        15'b111110011111010 : reciprocal = 1111111111111111;
        15'b111110011111001 : reciprocal = 1111111111111111;
        15'b111110011111000 : reciprocal = 1111111111111111;
        15'b111110011110111 : reciprocal = 1111111111111111;
        15'b111110011110110 : reciprocal = 1111111111111111;
        15'b111110011110101 : reciprocal = 1111111111111111;
        15'b111110011110100 : reciprocal = 1111111111111111;
        15'b111110011110011 : reciprocal = 1111111111111111;
        15'b111110011110010 : reciprocal = 1111111111111111;
        15'b111110011110001 : reciprocal = 1111111111111111;
        15'b111110011110000 : reciprocal = 1111111111111111;
        15'b111110011101111 : reciprocal = 1111111111111111;
        15'b111110011101110 : reciprocal = 1111111111111111;
        15'b111110011101101 : reciprocal = 1111111111111111;
        15'b111110011101100 : reciprocal = 1111111111111111;
        15'b111110011101011 : reciprocal = 1111111111111111;
        15'b111110011101010 : reciprocal = 1111111111111111;
        15'b111110011101001 : reciprocal = 1111111111111111;
        15'b111110011101000 : reciprocal = 1111111111111111;
        15'b111110011100111 : reciprocal = 1111111111111111;
        15'b111110011100110 : reciprocal = 1111111111111111;
        15'b111110011100101 : reciprocal = 1111111111111111;
        15'b111110011100100 : reciprocal = 1111111111111111;
        15'b111110011100011 : reciprocal = 1111111111111111;
        15'b111110011100010 : reciprocal = 1111111111111111;
        15'b111110011100001 : reciprocal = 1111111111111111;
        15'b111110011100000 : reciprocal = 1111111111111111;
        15'b111110011011111 : reciprocal = 1111111111111111;
        15'b111110011011110 : reciprocal = 1111111111111111;
        15'b111110011011101 : reciprocal = 1111111111111111;
        15'b111110011011100 : reciprocal = 1111111111111111;
        15'b111110011011011 : reciprocal = 1111111111111111;
        15'b111110011011010 : reciprocal = 1111111111111111;
        15'b111110011011001 : reciprocal = 1111111111111111;
        15'b111110011011000 : reciprocal = 1111111111111111;
        15'b111110011010111 : reciprocal = 1111111111111111;
        15'b111110011010110 : reciprocal = 1111111111111111;
        15'b111110011010101 : reciprocal = 1111111111111111;
        15'b111110011010100 : reciprocal = 1111111111111111;
        15'b111110011010011 : reciprocal = 1111111111111111;
        15'b111110011010010 : reciprocal = 1111111111111111;
        15'b111110011010001 : reciprocal = 1111111111111111;
        15'b111110011010000 : reciprocal = 1111111111111111;
        15'b111110011001111 : reciprocal = 1111111111111111;
        15'b111110011001110 : reciprocal = 1111111111111111;
        15'b111110011001101 : reciprocal = 1111111111111111;
        15'b111110011001100 : reciprocal = 1111111111111111;
        15'b111110011001011 : reciprocal = 1111111111111111;
        15'b111110011001010 : reciprocal = 1111111111111111;
        15'b111110011001001 : reciprocal = 1111111111111111;
        15'b111110011001000 : reciprocal = 1111111111111111;
        15'b111110011000111 : reciprocal = 1111111111111111;
        15'b111110011000110 : reciprocal = 1111111111111111;
        15'b111110011000101 : reciprocal = 1111111111111111;
        15'b111110011000100 : reciprocal = 1111111111111111;
        15'b111110011000011 : reciprocal = 1111111111111111;
        15'b111110011000010 : reciprocal = 1111111111111111;
        15'b111110011000001 : reciprocal = 1111111111111111;
        15'b111110011000000 : reciprocal = 1111111111111111;
        15'b111110010111111 : reciprocal = 1111111111111111;
        15'b111110010111110 : reciprocal = 1111111111111111;
        15'b111110010111101 : reciprocal = 1111111111111111;
        15'b111110010111100 : reciprocal = 1111111111111111;
        15'b111110010111011 : reciprocal = 1111111111111111;
        15'b111110010111010 : reciprocal = 1111111111111111;
        15'b111110010111001 : reciprocal = 1111111111111111;
        15'b111110010111000 : reciprocal = 1111111111111111;
        15'b111110010110111 : reciprocal = 1111111111111111;
        15'b111110010110110 : reciprocal = 1111111111111111;
        15'b111110010110101 : reciprocal = 1111111111111111;
        15'b111110010110100 : reciprocal = 1111111111111111;
        15'b111110010110011 : reciprocal = 1111111111111111;
        15'b111110010110010 : reciprocal = 1111111111111111;
        15'b111110010110001 : reciprocal = 1111111111111111;
        15'b111110010110000 : reciprocal = 1111111111111111;
        15'b111110010101111 : reciprocal = 1111111111111111;
        15'b111110010101110 : reciprocal = 1111111111111111;
        15'b111110010101101 : reciprocal = 1111111111111111;
        15'b111110010101100 : reciprocal = 1111111111111111;
        15'b111110010101011 : reciprocal = 1111111111111111;
        15'b111110010101010 : reciprocal = 1111111111111111;
        15'b111110010101001 : reciprocal = 1111111111111111;
        15'b111110010101000 : reciprocal = 1111111111111111;
        15'b111110010100111 : reciprocal = 1111111111111111;
        15'b111110010100110 : reciprocal = 1111111111111111;
        15'b111110010100101 : reciprocal = 1111111111111111;
        15'b111110010100100 : reciprocal = 1111111111111111;
        15'b111110010100011 : reciprocal = 1111111111111111;
        15'b111110010100010 : reciprocal = 1111111111111111;
        15'b111110010100001 : reciprocal = 1111111111111111;
        15'b111110010100000 : reciprocal = 1111111111111111;
        15'b111110010011111 : reciprocal = 1111111111111111;
        15'b111110010011110 : reciprocal = 1111111111111111;
        15'b111110010011101 : reciprocal = 1111111111111111;
        15'b111110010011100 : reciprocal = 1111111111111111;
        15'b111110010011011 : reciprocal = 1111111111111111;
        15'b111110010011010 : reciprocal = 1111111111111111;
        15'b111110010011001 : reciprocal = 1111111111111111;
        15'b111110010011000 : reciprocal = 1111111111111111;
        15'b111110010010111 : reciprocal = 1111111111111111;
        15'b111110010010110 : reciprocal = 1111111111111111;
        15'b111110010010101 : reciprocal = 1111111111111111;
        15'b111110010010100 : reciprocal = 1111111111111111;
        15'b111110010010011 : reciprocal = 1111111111111111;
        15'b111110010010010 : reciprocal = 1111111111111111;
        15'b111110010010001 : reciprocal = 1111111111111111;
        15'b111110010010000 : reciprocal = 1111111111111111;
        15'b111110010001111 : reciprocal = 1111111111111111;
        15'b111110010001110 : reciprocal = 1111111111111111;
        15'b111110010001101 : reciprocal = 1111111111111111;
        15'b111110010001100 : reciprocal = 1111111111111111;
        15'b111110010001011 : reciprocal = 1111111111111111;
        15'b111110010001010 : reciprocal = 1111111111111111;
        15'b111110010001001 : reciprocal = 1111111111111111;
        15'b111110010001000 : reciprocal = 1111111111111111;
        15'b111110010000111 : reciprocal = 1111111111111111;
        15'b111110010000110 : reciprocal = 1111111111111111;
        15'b111110010000101 : reciprocal = 1111111111111111;
        15'b111110010000100 : reciprocal = 1111111111111111;
        15'b111110010000011 : reciprocal = 1111111111111111;
        15'b111110010000010 : reciprocal = 1111111111111111;
        15'b111110010000001 : reciprocal = 1111111111111111;
        15'b111110010000000 : reciprocal = 1111111111111111;
        15'b111110001111111 : reciprocal = 1111111111111111;
        15'b111110001111110 : reciprocal = 1111111111111111;
        15'b111110001111101 : reciprocal = 1111111111111111;
        15'b111110001111100 : reciprocal = 1111111111111111;
        15'b111110001111011 : reciprocal = 1111111111111111;
        15'b111110001111010 : reciprocal = 1111111111111111;
        15'b111110001111001 : reciprocal = 1111111111111111;
        15'b111110001111000 : reciprocal = 1111111111111111;
        15'b111110001110111 : reciprocal = 1111111111111111;
        15'b111110001110110 : reciprocal = 1111111111111111;
        15'b111110001110101 : reciprocal = 1111111111111111;
        15'b111110001110100 : reciprocal = 1111111111111111;
        15'b111110001110011 : reciprocal = 1111111111111111;
        15'b111110001110010 : reciprocal = 1111111111111111;
        15'b111110001110001 : reciprocal = 1111111111111111;
        15'b111110001110000 : reciprocal = 1111111111111111;
        15'b111110001101111 : reciprocal = 1111111111111111;
        15'b111110001101110 : reciprocal = 1111111111111111;
        15'b111110001101101 : reciprocal = 1111111111111111;
        15'b111110001101100 : reciprocal = 1111111111111111;
        15'b111110001101011 : reciprocal = 1111111111111111;
        15'b111110001101010 : reciprocal = 1111111111111111;
        15'b111110001101001 : reciprocal = 1111111111111111;
        15'b111110001101000 : reciprocal = 1111111111111111;
        15'b111110001100111 : reciprocal = 1111111111111111;
        15'b111110001100110 : reciprocal = 1111111111111111;
        15'b111110001100101 : reciprocal = 1111111111111111;
        15'b111110001100100 : reciprocal = 1111111111111111;
        15'b111110001100011 : reciprocal = 1111111111111111;
        15'b111110001100010 : reciprocal = 1111111111111111;
        15'b111110001100001 : reciprocal = 1111111111111111;
        15'b111110001100000 : reciprocal = 1111111111111111;
        15'b111110001011111 : reciprocal = 1111111111111111;
        15'b111110001011110 : reciprocal = 1111111111111111;
        15'b111110001011101 : reciprocal = 1111111111111111;
        15'b111110001011100 : reciprocal = 1111111111111111;
        15'b111110001011011 : reciprocal = 1111111111111111;
        15'b111110001011010 : reciprocal = 1111111111111111;
        15'b111110001011001 : reciprocal = 1111111111111111;
        15'b111110001011000 : reciprocal = 1111111111111111;
        15'b111110001010111 : reciprocal = 1111111111111111;
        15'b111110001010110 : reciprocal = 1111111111111111;
        15'b111110001010101 : reciprocal = 1111111111111111;
        15'b111110001010100 : reciprocal = 1111111111111111;
        15'b111110001010011 : reciprocal = 1111111111111111;
        15'b111110001010010 : reciprocal = 1111111111111111;
        15'b111110001010001 : reciprocal = 1111111111111111;
        15'b111110001010000 : reciprocal = 1111111111111111;
        15'b111110001001111 : reciprocal = 1111111111111111;
        15'b111110001001110 : reciprocal = 1111111111111111;
        15'b111110001001101 : reciprocal = 1111111111111111;
        15'b111110001001100 : reciprocal = 1111111111111111;
        15'b111110001001011 : reciprocal = 1111111111111111;
        15'b111110001001010 : reciprocal = 1111111111111111;
        15'b111110001001001 : reciprocal = 1111111111111111;
        15'b111110001001000 : reciprocal = 1111111111111111;
        15'b111110001000111 : reciprocal = 1111111111111111;
        15'b111110001000110 : reciprocal = 1111111111111111;
        15'b111110001000101 : reciprocal = 1111111111111111;
        15'b111110001000100 : reciprocal = 1111111111111111;
        15'b111110001000011 : reciprocal = 1111111111111111;
        15'b111110001000010 : reciprocal = 1111111111111111;
        15'b111110001000001 : reciprocal = 1111111111111111;
        15'b111110001000000 : reciprocal = 1111111111111111;
        15'b111110000111111 : reciprocal = 1111111111111111;
        15'b111110000111110 : reciprocal = 1111111111111111;
        15'b111110000111101 : reciprocal = 1111111111111111;
        15'b111110000111100 : reciprocal = 1111111111111111;
        15'b111110000111011 : reciprocal = 1111111111111111;
        15'b111110000111010 : reciprocal = 1111111111111111;
        15'b111110000111001 : reciprocal = 1111111111111111;
        15'b111110000111000 : reciprocal = 1111111111111111;
        15'b111110000110111 : reciprocal = 1111111111111111;
        15'b111110000110110 : reciprocal = 1111111111111111;
        15'b111110000110101 : reciprocal = 1111111111111111;
        15'b111110000110100 : reciprocal = 1111111111111111;
        15'b111110000110011 : reciprocal = 1111111111111111;
        15'b111110000110010 : reciprocal = 1111111111111111;
        15'b111110000110001 : reciprocal = 1111111111111111;
        15'b111110000110000 : reciprocal = 1111111111111111;
        15'b111110000101111 : reciprocal = 1111111111111111;
        15'b111110000101110 : reciprocal = 1111111111111111;
        15'b111110000101101 : reciprocal = 1111111111111111;
        15'b111110000101100 : reciprocal = 1111111111111111;
        15'b111110000101011 : reciprocal = 1111111111111111;
        15'b111110000101010 : reciprocal = 1111111111111111;
        15'b111110000101001 : reciprocal = 1111111111111111;
        15'b111110000101000 : reciprocal = 1111111111111111;
        15'b111110000100111 : reciprocal = 1111111111111111;
        15'b111110000100110 : reciprocal = 1111111111111111;
        15'b111110000100101 : reciprocal = 1111111111111111;
        15'b111110000100100 : reciprocal = 1111111111111111;
        15'b111110000100011 : reciprocal = 1111111111111111;
        15'b111110000100010 : reciprocal = 1111111111111111;
        15'b111110000100001 : reciprocal = 1111111111111111;
        15'b111110000100000 : reciprocal = 1111111111111111;
        15'b111110000011111 : reciprocal = 1111111111111111;
        15'b111110000011110 : reciprocal = 1111111111111111;
        15'b111110000011101 : reciprocal = 1111111111111111;
        15'b111110000011100 : reciprocal = 1111111111111111;
        15'b111110000011011 : reciprocal = 1111111111111111;
        15'b111110000011010 : reciprocal = 1111111111111111;
        15'b111110000011001 : reciprocal = 1111111111111111;
        15'b111110000011000 : reciprocal = 1111111111111111;
        15'b111110000010111 : reciprocal = 1111111111111111;
        15'b111110000010110 : reciprocal = 1111111111111111;
        15'b111110000010101 : reciprocal = 1111111111111111;
        15'b111110000010100 : reciprocal = 1111111111111111;
        15'b111110000010011 : reciprocal = 1111111111111111;
        15'b111110000010010 : reciprocal = 1111111111111111;
        15'b111110000010001 : reciprocal = 1111111111111111;
        15'b111110000010000 : reciprocal = 1111111111111111;
        15'b111110000001111 : reciprocal = 1111111111111111;
        15'b111110000001110 : reciprocal = 1111111111111111;
        15'b111110000001101 : reciprocal = 1111111111111111;
        15'b111110000001100 : reciprocal = 1111111111111111;
        15'b111110000001011 : reciprocal = 1111111111111111;
        15'b111110000001010 : reciprocal = 1111111111111111;
        15'b111110000001001 : reciprocal = 1111111111111111;
        15'b111110000001000 : reciprocal = 1111111111111111;
        15'b111110000000111 : reciprocal = 1111111111111111;
        15'b111110000000110 : reciprocal = 1111111111111111;
        15'b111110000000101 : reciprocal = 1111111111111111;
        15'b111110000000100 : reciprocal = 1111111111111111;
        15'b111110000000011 : reciprocal = 1111111111111111;
        15'b111110000000010 : reciprocal = 1111111111111111;
        15'b111110000000001 : reciprocal = 1111111111111111;


        endcase
    end
    



    //////////////////////// For testbenching ////////////////////////
    // synthesis translate_off

    // synthesis translate_on

endmodule
