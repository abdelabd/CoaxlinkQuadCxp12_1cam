module division_LUT_ap_fixed_16_10_s16 #(
)(
    input logic [16-1:0] number_in,
    output logic [16-1:0] reciprocal

);

    logic [65535:0] reciprocal_LUT [16-1:0];

    always_comb begin
        case (number_in[16-1:16-16])
        16'b0000000000000001 : reciprocal = 16'b0000010000000000;
        16'b0000000000000010 : reciprocal = 16'b0000001000000000;
        16'b0000000000000011 : reciprocal = 16'b0000000101010101;
        16'b0000000000000100 : reciprocal = 16'b0000000100000000;
        16'b0000000000000101 : reciprocal = 16'b0000000011001101;
        16'b0000000000000110 : reciprocal = 16'b0000000010101011;
        16'b0000000000000111 : reciprocal = 16'b0000000010010010;
        16'b0000000000001000 : reciprocal = 16'b0000000010000000;
        16'b0000000000001001 : reciprocal = 16'b0000000001110010;
        16'b0000000000001010 : reciprocal = 16'b0000000001100110;
        16'b0000000000001011 : reciprocal = 16'b0000000001011101;
        16'b0000000000001100 : reciprocal = 16'b0000000001010101;
        16'b0000000000001101 : reciprocal = 16'b0000000001001111;
        16'b0000000000001110 : reciprocal = 16'b0000000001001001;
        16'b0000000000001111 : reciprocal = 16'b0000000001000100;
        16'b0000000000010000 : reciprocal = 16'b0000000001000000;
        16'b0000000000010001 : reciprocal = 16'b0000000000111100;
        16'b0000000000010010 : reciprocal = 16'b0000000000111001;
        16'b0000000000010011 : reciprocal = 16'b0000000000110110;
        16'b0000000000010100 : reciprocal = 16'b0000000000110011;
        16'b0000000000010101 : reciprocal = 16'b0000000000110001;
        16'b0000000000010110 : reciprocal = 16'b0000000000101111;
        16'b0000000000010111 : reciprocal = 16'b0000000000101101;
        16'b0000000000011000 : reciprocal = 16'b0000000000101011;
        16'b0000000000011001 : reciprocal = 16'b0000000000101001;
        16'b0000000000011010 : reciprocal = 16'b0000000000100111;
        16'b0000000000011011 : reciprocal = 16'b0000000000100110;
        16'b0000000000011100 : reciprocal = 16'b0000000000100101;
        16'b0000000000011101 : reciprocal = 16'b0000000000100011;
        16'b0000000000011110 : reciprocal = 16'b0000000000100010;
        16'b0000000000011111 : reciprocal = 16'b0000000000100001;
        16'b0000000000100000 : reciprocal = 16'b0000000000100000;
        16'b0000000000100001 : reciprocal = 16'b0000000000011111;
        16'b0000000000100010 : reciprocal = 16'b0000000000011110;
        16'b0000000000100011 : reciprocal = 16'b0000000000011101;
        16'b0000000000100100 : reciprocal = 16'b0000000000011100;
        16'b0000000000100101 : reciprocal = 16'b0000000000011100;
        16'b0000000000100110 : reciprocal = 16'b0000000000011011;
        16'b0000000000100111 : reciprocal = 16'b0000000000011010;
        16'b0000000000101000 : reciprocal = 16'b0000000000011010;
        16'b0000000000101001 : reciprocal = 16'b0000000000011001;
        16'b0000000000101010 : reciprocal = 16'b0000000000011000;
        16'b0000000000101011 : reciprocal = 16'b0000000000011000;
        16'b0000000000101100 : reciprocal = 16'b0000000000010111;
        16'b0000000000101101 : reciprocal = 16'b0000000000010111;
        16'b0000000000101110 : reciprocal = 16'b0000000000010110;
        16'b0000000000101111 : reciprocal = 16'b0000000000010110;
        16'b0000000000110000 : reciprocal = 16'b0000000000010101;
        16'b0000000000110001 : reciprocal = 16'b0000000000010101;
        16'b0000000000110010 : reciprocal = 16'b0000000000010100;
        16'b0000000000110011 : reciprocal = 16'b0000000000010100;
        16'b0000000000110100 : reciprocal = 16'b0000000000010100;
        16'b0000000000110101 : reciprocal = 16'b0000000000010011;
        16'b0000000000110110 : reciprocal = 16'b0000000000010011;
        16'b0000000000110111 : reciprocal = 16'b0000000000010011;
        16'b0000000000111000 : reciprocal = 16'b0000000000010010;
        16'b0000000000111001 : reciprocal = 16'b0000000000010010;
        16'b0000000000111010 : reciprocal = 16'b0000000000010010;
        16'b0000000000111011 : reciprocal = 16'b0000000000010001;
        16'b0000000000111100 : reciprocal = 16'b0000000000010001;
        16'b0000000000111101 : reciprocal = 16'b0000000000010001;
        16'b0000000000111110 : reciprocal = 16'b0000000000010001;
        16'b0000000000111111 : reciprocal = 16'b0000000000010000;
        16'b0000000001000000 : reciprocal = 16'b0000000000010000;
        16'b0000000001000001 : reciprocal = 16'b0000000000010000;
        16'b0000000001000010 : reciprocal = 16'b0000000000010000;
        16'b0000000001000011 : reciprocal = 16'b0000000000001111;
        16'b0000000001000100 : reciprocal = 16'b0000000000001111;
        16'b0000000001000101 : reciprocal = 16'b0000000000001111;
        16'b0000000001000110 : reciprocal = 16'b0000000000001111;
        16'b0000000001000111 : reciprocal = 16'b0000000000001110;
        16'b0000000001001000 : reciprocal = 16'b0000000000001110;
        16'b0000000001001001 : reciprocal = 16'b0000000000001110;
        16'b0000000001001010 : reciprocal = 16'b0000000000001110;
        16'b0000000001001011 : reciprocal = 16'b0000000000001110;
        16'b0000000001001100 : reciprocal = 16'b0000000000001101;
        16'b0000000001001101 : reciprocal = 16'b0000000000001101;
        16'b0000000001001110 : reciprocal = 16'b0000000000001101;
        16'b0000000001001111 : reciprocal = 16'b0000000000001101;
        16'b0000000001010000 : reciprocal = 16'b0000000000001101;
        16'b0000000001010001 : reciprocal = 16'b0000000000001101;
        16'b0000000001010010 : reciprocal = 16'b0000000000001100;
        16'b0000000001010011 : reciprocal = 16'b0000000000001100;
        16'b0000000001010100 : reciprocal = 16'b0000000000001100;
        16'b0000000001010101 : reciprocal = 16'b0000000000001100;
        16'b0000000001010110 : reciprocal = 16'b0000000000001100;
        16'b0000000001010111 : reciprocal = 16'b0000000000001100;
        16'b0000000001011000 : reciprocal = 16'b0000000000001100;
        16'b0000000001011001 : reciprocal = 16'b0000000000001100;
        16'b0000000001011010 : reciprocal = 16'b0000000000001011;
        16'b0000000001011011 : reciprocal = 16'b0000000000001011;
        16'b0000000001011100 : reciprocal = 16'b0000000000001011;
        16'b0000000001011101 : reciprocal = 16'b0000000000001011;
        16'b0000000001011110 : reciprocal = 16'b0000000000001011;
        16'b0000000001011111 : reciprocal = 16'b0000000000001011;
        16'b0000000001100000 : reciprocal = 16'b0000000000001011;
        16'b0000000001100001 : reciprocal = 16'b0000000000001011;
        16'b0000000001100010 : reciprocal = 16'b0000000000001010;
        16'b0000000001100011 : reciprocal = 16'b0000000000001010;
        16'b0000000001100100 : reciprocal = 16'b0000000000001010;
        16'b0000000001100101 : reciprocal = 16'b0000000000001010;
        16'b0000000001100110 : reciprocal = 16'b0000000000001010;
        16'b0000000001100111 : reciprocal = 16'b0000000000001010;
        16'b0000000001101000 : reciprocal = 16'b0000000000001010;
        16'b0000000001101001 : reciprocal = 16'b0000000000001010;
        16'b0000000001101010 : reciprocal = 16'b0000000000001010;
        16'b0000000001101011 : reciprocal = 16'b0000000000001010;
        16'b0000000001101100 : reciprocal = 16'b0000000000001001;
        16'b0000000001101101 : reciprocal = 16'b0000000000001001;
        16'b0000000001101110 : reciprocal = 16'b0000000000001001;
        16'b0000000001101111 : reciprocal = 16'b0000000000001001;
        16'b0000000001110000 : reciprocal = 16'b0000000000001001;
        16'b0000000001110001 : reciprocal = 16'b0000000000001001;
        16'b0000000001110010 : reciprocal = 16'b0000000000001001;
        16'b0000000001110011 : reciprocal = 16'b0000000000001001;
        16'b0000000001110100 : reciprocal = 16'b0000000000001001;
        16'b0000000001110101 : reciprocal = 16'b0000000000001001;
        16'b0000000001110110 : reciprocal = 16'b0000000000001001;
        16'b0000000001110111 : reciprocal = 16'b0000000000001001;
        16'b0000000001111000 : reciprocal = 16'b0000000000001001;
        16'b0000000001111001 : reciprocal = 16'b0000000000001000;
        16'b0000000001111010 : reciprocal = 16'b0000000000001000;
        16'b0000000001111011 : reciprocal = 16'b0000000000001000;
        16'b0000000001111100 : reciprocal = 16'b0000000000001000;
        16'b0000000001111101 : reciprocal = 16'b0000000000001000;
        16'b0000000001111110 : reciprocal = 16'b0000000000001000;
        16'b0000000001111111 : reciprocal = 16'b0000000000001000;
        16'b0000000010000000 : reciprocal = 16'b0000000000001000;
        16'b0000000010000001 : reciprocal = 16'b0000000000001000;
        16'b0000000010000010 : reciprocal = 16'b0000000000001000;
        16'b0000000010000011 : reciprocal = 16'b0000000000001000;
        16'b0000000010000100 : reciprocal = 16'b0000000000001000;
        16'b0000000010000101 : reciprocal = 16'b0000000000001000;
        16'b0000000010000110 : reciprocal = 16'b0000000000001000;
        16'b0000000010000111 : reciprocal = 16'b0000000000001000;
        16'b0000000010001000 : reciprocal = 16'b0000000000001000;
        16'b0000000010001001 : reciprocal = 16'b0000000000000111;
        16'b0000000010001010 : reciprocal = 16'b0000000000000111;
        16'b0000000010001011 : reciprocal = 16'b0000000000000111;
        16'b0000000010001100 : reciprocal = 16'b0000000000000111;
        16'b0000000010001101 : reciprocal = 16'b0000000000000111;
        16'b0000000010001110 : reciprocal = 16'b0000000000000111;
        16'b0000000010001111 : reciprocal = 16'b0000000000000111;
        16'b0000000010010000 : reciprocal = 16'b0000000000000111;
        16'b0000000010010001 : reciprocal = 16'b0000000000000111;
        16'b0000000010010010 : reciprocal = 16'b0000000000000111;
        16'b0000000010010011 : reciprocal = 16'b0000000000000111;
        16'b0000000010010100 : reciprocal = 16'b0000000000000111;
        16'b0000000010010101 : reciprocal = 16'b0000000000000111;
        16'b0000000010010110 : reciprocal = 16'b0000000000000111;
        16'b0000000010010111 : reciprocal = 16'b0000000000000111;
        16'b0000000010011000 : reciprocal = 16'b0000000000000111;
        16'b0000000010011001 : reciprocal = 16'b0000000000000111;
        16'b0000000010011010 : reciprocal = 16'b0000000000000111;
        16'b0000000010011011 : reciprocal = 16'b0000000000000111;
        16'b0000000010011100 : reciprocal = 16'b0000000000000111;
        16'b0000000010011101 : reciprocal = 16'b0000000000000111;
        16'b0000000010011110 : reciprocal = 16'b0000000000000110;
        16'b0000000010011111 : reciprocal = 16'b0000000000000110;
        16'b0000000010100000 : reciprocal = 16'b0000000000000110;
        16'b0000000010100001 : reciprocal = 16'b0000000000000110;
        16'b0000000010100010 : reciprocal = 16'b0000000000000110;
        16'b0000000010100011 : reciprocal = 16'b0000000000000110;
        16'b0000000010100100 : reciprocal = 16'b0000000000000110;
        16'b0000000010100101 : reciprocal = 16'b0000000000000110;
        16'b0000000010100110 : reciprocal = 16'b0000000000000110;
        16'b0000000010100111 : reciprocal = 16'b0000000000000110;
        16'b0000000010101000 : reciprocal = 16'b0000000000000110;
        16'b0000000010101001 : reciprocal = 16'b0000000000000110;
        16'b0000000010101010 : reciprocal = 16'b0000000000000110;
        16'b0000000010101011 : reciprocal = 16'b0000000000000110;
        16'b0000000010101100 : reciprocal = 16'b0000000000000110;
        16'b0000000010101101 : reciprocal = 16'b0000000000000110;
        16'b0000000010101110 : reciprocal = 16'b0000000000000110;
        16'b0000000010101111 : reciprocal = 16'b0000000000000110;
        16'b0000000010110000 : reciprocal = 16'b0000000000000110;
        16'b0000000010110001 : reciprocal = 16'b0000000000000110;
        16'b0000000010110010 : reciprocal = 16'b0000000000000110;
        16'b0000000010110011 : reciprocal = 16'b0000000000000110;
        16'b0000000010110100 : reciprocal = 16'b0000000000000110;
        16'b0000000010110101 : reciprocal = 16'b0000000000000110;
        16'b0000000010110110 : reciprocal = 16'b0000000000000110;
        16'b0000000010110111 : reciprocal = 16'b0000000000000110;
        16'b0000000010111000 : reciprocal = 16'b0000000000000110;
        16'b0000000010111001 : reciprocal = 16'b0000000000000110;
        16'b0000000010111010 : reciprocal = 16'b0000000000000110;
        16'b0000000010111011 : reciprocal = 16'b0000000000000101;
        16'b0000000010111100 : reciprocal = 16'b0000000000000101;
        16'b0000000010111101 : reciprocal = 16'b0000000000000101;
        16'b0000000010111110 : reciprocal = 16'b0000000000000101;
        16'b0000000010111111 : reciprocal = 16'b0000000000000101;
        16'b0000000011000000 : reciprocal = 16'b0000000000000101;
        16'b0000000011000001 : reciprocal = 16'b0000000000000101;
        16'b0000000011000010 : reciprocal = 16'b0000000000000101;
        16'b0000000011000011 : reciprocal = 16'b0000000000000101;
        16'b0000000011000100 : reciprocal = 16'b0000000000000101;
        16'b0000000011000101 : reciprocal = 16'b0000000000000101;
        16'b0000000011000110 : reciprocal = 16'b0000000000000101;
        16'b0000000011000111 : reciprocal = 16'b0000000000000101;
        16'b0000000011001000 : reciprocal = 16'b0000000000000101;
        16'b0000000011001001 : reciprocal = 16'b0000000000000101;
        16'b0000000011001010 : reciprocal = 16'b0000000000000101;
        16'b0000000011001011 : reciprocal = 16'b0000000000000101;
        16'b0000000011001100 : reciprocal = 16'b0000000000000101;
        16'b0000000011001101 : reciprocal = 16'b0000000000000101;
        16'b0000000011001110 : reciprocal = 16'b0000000000000101;
        16'b0000000011001111 : reciprocal = 16'b0000000000000101;
        16'b0000000011010000 : reciprocal = 16'b0000000000000101;
        16'b0000000011010001 : reciprocal = 16'b0000000000000101;
        16'b0000000011010010 : reciprocal = 16'b0000000000000101;
        16'b0000000011010011 : reciprocal = 16'b0000000000000101;
        16'b0000000011010100 : reciprocal = 16'b0000000000000101;
        16'b0000000011010101 : reciprocal = 16'b0000000000000101;
        16'b0000000011010110 : reciprocal = 16'b0000000000000101;
        16'b0000000011010111 : reciprocal = 16'b0000000000000101;
        16'b0000000011011000 : reciprocal = 16'b0000000000000101;
        16'b0000000011011001 : reciprocal = 16'b0000000000000101;
        16'b0000000011011010 : reciprocal = 16'b0000000000000101;
        16'b0000000011011011 : reciprocal = 16'b0000000000000101;
        16'b0000000011011100 : reciprocal = 16'b0000000000000101;
        16'b0000000011011101 : reciprocal = 16'b0000000000000101;
        16'b0000000011011110 : reciprocal = 16'b0000000000000101;
        16'b0000000011011111 : reciprocal = 16'b0000000000000101;
        16'b0000000011100000 : reciprocal = 16'b0000000000000101;
        16'b0000000011100001 : reciprocal = 16'b0000000000000101;
        16'b0000000011100010 : reciprocal = 16'b0000000000000101;
        16'b0000000011100011 : reciprocal = 16'b0000000000000101;
        16'b0000000011100100 : reciprocal = 16'b0000000000000100;
        16'b0000000011100101 : reciprocal = 16'b0000000000000100;
        16'b0000000011100110 : reciprocal = 16'b0000000000000100;
        16'b0000000011100111 : reciprocal = 16'b0000000000000100;
        16'b0000000011101000 : reciprocal = 16'b0000000000000100;
        16'b0000000011101001 : reciprocal = 16'b0000000000000100;
        16'b0000000011101010 : reciprocal = 16'b0000000000000100;
        16'b0000000011101011 : reciprocal = 16'b0000000000000100;
        16'b0000000011101100 : reciprocal = 16'b0000000000000100;
        16'b0000000011101101 : reciprocal = 16'b0000000000000100;
        16'b0000000011101110 : reciprocal = 16'b0000000000000100;
        16'b0000000011101111 : reciprocal = 16'b0000000000000100;
        16'b0000000011110000 : reciprocal = 16'b0000000000000100;
        16'b0000000011110001 : reciprocal = 16'b0000000000000100;
        16'b0000000011110010 : reciprocal = 16'b0000000000000100;
        16'b0000000011110011 : reciprocal = 16'b0000000000000100;
        16'b0000000011110100 : reciprocal = 16'b0000000000000100;
        16'b0000000011110101 : reciprocal = 16'b0000000000000100;
        16'b0000000011110110 : reciprocal = 16'b0000000000000100;
        16'b0000000011110111 : reciprocal = 16'b0000000000000100;
        16'b0000000011111000 : reciprocal = 16'b0000000000000100;
        16'b0000000011111001 : reciprocal = 16'b0000000000000100;
        16'b0000000011111010 : reciprocal = 16'b0000000000000100;
        16'b0000000011111011 : reciprocal = 16'b0000000000000100;
        16'b0000000011111100 : reciprocal = 16'b0000000000000100;
        16'b0000000011111101 : reciprocal = 16'b0000000000000100;
        16'b0000000011111110 : reciprocal = 16'b0000000000000100;
        16'b0000000011111111 : reciprocal = 16'b0000000000000100;
        16'b0000000100000000 : reciprocal = 16'b0000000000000100;
        16'b0000000100000001 : reciprocal = 16'b0000000000000100;
        16'b0000000100000010 : reciprocal = 16'b0000000000000100;
        16'b0000000100000011 : reciprocal = 16'b0000000000000100;
        16'b0000000100000100 : reciprocal = 16'b0000000000000100;
        16'b0000000100000101 : reciprocal = 16'b0000000000000100;
        16'b0000000100000110 : reciprocal = 16'b0000000000000100;
        16'b0000000100000111 : reciprocal = 16'b0000000000000100;
        16'b0000000100001000 : reciprocal = 16'b0000000000000100;
        16'b0000000100001001 : reciprocal = 16'b0000000000000100;
        16'b0000000100001010 : reciprocal = 16'b0000000000000100;
        16'b0000000100001011 : reciprocal = 16'b0000000000000100;
        16'b0000000100001100 : reciprocal = 16'b0000000000000100;
        16'b0000000100001101 : reciprocal = 16'b0000000000000100;
        16'b0000000100001110 : reciprocal = 16'b0000000000000100;
        16'b0000000100001111 : reciprocal = 16'b0000000000000100;
        16'b0000000100010000 : reciprocal = 16'b0000000000000100;
        16'b0000000100010001 : reciprocal = 16'b0000000000000100;
        16'b0000000100010010 : reciprocal = 16'b0000000000000100;
        16'b0000000100010011 : reciprocal = 16'b0000000000000100;
        16'b0000000100010100 : reciprocal = 16'b0000000000000100;
        16'b0000000100010101 : reciprocal = 16'b0000000000000100;
        16'b0000000100010110 : reciprocal = 16'b0000000000000100;
        16'b0000000100010111 : reciprocal = 16'b0000000000000100;
        16'b0000000100011000 : reciprocal = 16'b0000000000000100;
        16'b0000000100011001 : reciprocal = 16'b0000000000000100;
        16'b0000000100011010 : reciprocal = 16'b0000000000000100;
        16'b0000000100011011 : reciprocal = 16'b0000000000000100;
        16'b0000000100011100 : reciprocal = 16'b0000000000000100;
        16'b0000000100011101 : reciprocal = 16'b0000000000000100;
        16'b0000000100011110 : reciprocal = 16'b0000000000000100;
        16'b0000000100011111 : reciprocal = 16'b0000000000000100;
        16'b0000000100100000 : reciprocal = 16'b0000000000000100;
        16'b0000000100100001 : reciprocal = 16'b0000000000000100;
        16'b0000000100100010 : reciprocal = 16'b0000000000000100;
        16'b0000000100100011 : reciprocal = 16'b0000000000000100;
        16'b0000000100100100 : reciprocal = 16'b0000000000000100;
        16'b0000000100100101 : reciprocal = 16'b0000000000000011;
        16'b0000000100100110 : reciprocal = 16'b0000000000000011;
        16'b0000000100100111 : reciprocal = 16'b0000000000000011;
        16'b0000000100101000 : reciprocal = 16'b0000000000000011;
        16'b0000000100101001 : reciprocal = 16'b0000000000000011;
        16'b0000000100101010 : reciprocal = 16'b0000000000000011;
        16'b0000000100101011 : reciprocal = 16'b0000000000000011;
        16'b0000000100101100 : reciprocal = 16'b0000000000000011;
        16'b0000000100101101 : reciprocal = 16'b0000000000000011;
        16'b0000000100101110 : reciprocal = 16'b0000000000000011;
        16'b0000000100101111 : reciprocal = 16'b0000000000000011;
        16'b0000000100110000 : reciprocal = 16'b0000000000000011;
        16'b0000000100110001 : reciprocal = 16'b0000000000000011;
        16'b0000000100110010 : reciprocal = 16'b0000000000000011;
        16'b0000000100110011 : reciprocal = 16'b0000000000000011;
        16'b0000000100110100 : reciprocal = 16'b0000000000000011;
        16'b0000000100110101 : reciprocal = 16'b0000000000000011;
        16'b0000000100110110 : reciprocal = 16'b0000000000000011;
        16'b0000000100110111 : reciprocal = 16'b0000000000000011;
        16'b0000000100111000 : reciprocal = 16'b0000000000000011;
        16'b0000000100111001 : reciprocal = 16'b0000000000000011;
        16'b0000000100111010 : reciprocal = 16'b0000000000000011;
        16'b0000000100111011 : reciprocal = 16'b0000000000000011;
        16'b0000000100111100 : reciprocal = 16'b0000000000000011;
        16'b0000000100111101 : reciprocal = 16'b0000000000000011;
        16'b0000000100111110 : reciprocal = 16'b0000000000000011;
        16'b0000000100111111 : reciprocal = 16'b0000000000000011;
        16'b0000000101000000 : reciprocal = 16'b0000000000000011;
        16'b0000000101000001 : reciprocal = 16'b0000000000000011;
        16'b0000000101000010 : reciprocal = 16'b0000000000000011;
        16'b0000000101000011 : reciprocal = 16'b0000000000000011;
        16'b0000000101000100 : reciprocal = 16'b0000000000000011;
        16'b0000000101000101 : reciprocal = 16'b0000000000000011;
        16'b0000000101000110 : reciprocal = 16'b0000000000000011;
        16'b0000000101000111 : reciprocal = 16'b0000000000000011;
        16'b0000000101001000 : reciprocal = 16'b0000000000000011;
        16'b0000000101001001 : reciprocal = 16'b0000000000000011;
        16'b0000000101001010 : reciprocal = 16'b0000000000000011;
        16'b0000000101001011 : reciprocal = 16'b0000000000000011;
        16'b0000000101001100 : reciprocal = 16'b0000000000000011;
        16'b0000000101001101 : reciprocal = 16'b0000000000000011;
        16'b0000000101001110 : reciprocal = 16'b0000000000000011;
        16'b0000000101001111 : reciprocal = 16'b0000000000000011;
        16'b0000000101010000 : reciprocal = 16'b0000000000000011;
        16'b0000000101010001 : reciprocal = 16'b0000000000000011;
        16'b0000000101010010 : reciprocal = 16'b0000000000000011;
        16'b0000000101010011 : reciprocal = 16'b0000000000000011;
        16'b0000000101010100 : reciprocal = 16'b0000000000000011;
        16'b0000000101010101 : reciprocal = 16'b0000000000000011;
        16'b0000000101010110 : reciprocal = 16'b0000000000000011;
        16'b0000000101010111 : reciprocal = 16'b0000000000000011;
        16'b0000000101011000 : reciprocal = 16'b0000000000000011;
        16'b0000000101011001 : reciprocal = 16'b0000000000000011;
        16'b0000000101011010 : reciprocal = 16'b0000000000000011;
        16'b0000000101011011 : reciprocal = 16'b0000000000000011;
        16'b0000000101011100 : reciprocal = 16'b0000000000000011;
        16'b0000000101011101 : reciprocal = 16'b0000000000000011;
        16'b0000000101011110 : reciprocal = 16'b0000000000000011;
        16'b0000000101011111 : reciprocal = 16'b0000000000000011;
        16'b0000000101100000 : reciprocal = 16'b0000000000000011;
        16'b0000000101100001 : reciprocal = 16'b0000000000000011;
        16'b0000000101100010 : reciprocal = 16'b0000000000000011;
        16'b0000000101100011 : reciprocal = 16'b0000000000000011;
        16'b0000000101100100 : reciprocal = 16'b0000000000000011;
        16'b0000000101100101 : reciprocal = 16'b0000000000000011;
        16'b0000000101100110 : reciprocal = 16'b0000000000000011;
        16'b0000000101100111 : reciprocal = 16'b0000000000000011;
        16'b0000000101101000 : reciprocal = 16'b0000000000000011;
        16'b0000000101101001 : reciprocal = 16'b0000000000000011;
        16'b0000000101101010 : reciprocal = 16'b0000000000000011;
        16'b0000000101101011 : reciprocal = 16'b0000000000000011;
        16'b0000000101101100 : reciprocal = 16'b0000000000000011;
        16'b0000000101101101 : reciprocal = 16'b0000000000000011;
        16'b0000000101101110 : reciprocal = 16'b0000000000000011;
        16'b0000000101101111 : reciprocal = 16'b0000000000000011;
        16'b0000000101110000 : reciprocal = 16'b0000000000000011;
        16'b0000000101110001 : reciprocal = 16'b0000000000000011;
        16'b0000000101110010 : reciprocal = 16'b0000000000000011;
        16'b0000000101110011 : reciprocal = 16'b0000000000000011;
        16'b0000000101110100 : reciprocal = 16'b0000000000000011;
        16'b0000000101110101 : reciprocal = 16'b0000000000000011;
        16'b0000000101110110 : reciprocal = 16'b0000000000000011;
        16'b0000000101110111 : reciprocal = 16'b0000000000000011;
        16'b0000000101111000 : reciprocal = 16'b0000000000000011;
        16'b0000000101111001 : reciprocal = 16'b0000000000000011;
        16'b0000000101111010 : reciprocal = 16'b0000000000000011;
        16'b0000000101111011 : reciprocal = 16'b0000000000000011;
        16'b0000000101111100 : reciprocal = 16'b0000000000000011;
        16'b0000000101111101 : reciprocal = 16'b0000000000000011;
        16'b0000000101111110 : reciprocal = 16'b0000000000000011;
        16'b0000000101111111 : reciprocal = 16'b0000000000000011;
        16'b0000000110000000 : reciprocal = 16'b0000000000000011;
        16'b0000000110000001 : reciprocal = 16'b0000000000000011;
        16'b0000000110000010 : reciprocal = 16'b0000000000000011;
        16'b0000000110000011 : reciprocal = 16'b0000000000000011;
        16'b0000000110000100 : reciprocal = 16'b0000000000000011;
        16'b0000000110000101 : reciprocal = 16'b0000000000000011;
        16'b0000000110000110 : reciprocal = 16'b0000000000000011;
        16'b0000000110000111 : reciprocal = 16'b0000000000000011;
        16'b0000000110001000 : reciprocal = 16'b0000000000000011;
        16'b0000000110001001 : reciprocal = 16'b0000000000000011;
        16'b0000000110001010 : reciprocal = 16'b0000000000000011;
        16'b0000000110001011 : reciprocal = 16'b0000000000000011;
        16'b0000000110001100 : reciprocal = 16'b0000000000000011;
        16'b0000000110001101 : reciprocal = 16'b0000000000000011;
        16'b0000000110001110 : reciprocal = 16'b0000000000000011;
        16'b0000000110001111 : reciprocal = 16'b0000000000000011;
        16'b0000000110010000 : reciprocal = 16'b0000000000000011;
        16'b0000000110010001 : reciprocal = 16'b0000000000000011;
        16'b0000000110010010 : reciprocal = 16'b0000000000000011;
        16'b0000000110010011 : reciprocal = 16'b0000000000000011;
        16'b0000000110010100 : reciprocal = 16'b0000000000000011;
        16'b0000000110010101 : reciprocal = 16'b0000000000000011;
        16'b0000000110010110 : reciprocal = 16'b0000000000000011;
        16'b0000000110010111 : reciprocal = 16'b0000000000000011;
        16'b0000000110011000 : reciprocal = 16'b0000000000000011;
        16'b0000000110011001 : reciprocal = 16'b0000000000000011;
        16'b0000000110011010 : reciprocal = 16'b0000000000000010;
        16'b0000000110011011 : reciprocal = 16'b0000000000000010;
        16'b0000000110011100 : reciprocal = 16'b0000000000000010;
        16'b0000000110011101 : reciprocal = 16'b0000000000000010;
        16'b0000000110011110 : reciprocal = 16'b0000000000000010;
        16'b0000000110011111 : reciprocal = 16'b0000000000000010;
        16'b0000000110100000 : reciprocal = 16'b0000000000000010;
        16'b0000000110100001 : reciprocal = 16'b0000000000000010;
        16'b0000000110100010 : reciprocal = 16'b0000000000000010;
        16'b0000000110100011 : reciprocal = 16'b0000000000000010;
        16'b0000000110100100 : reciprocal = 16'b0000000000000010;
        16'b0000000110100101 : reciprocal = 16'b0000000000000010;
        16'b0000000110100110 : reciprocal = 16'b0000000000000010;
        16'b0000000110100111 : reciprocal = 16'b0000000000000010;
        16'b0000000110101000 : reciprocal = 16'b0000000000000010;
        16'b0000000110101001 : reciprocal = 16'b0000000000000010;
        16'b0000000110101010 : reciprocal = 16'b0000000000000010;
        16'b0000000110101011 : reciprocal = 16'b0000000000000010;
        16'b0000000110101100 : reciprocal = 16'b0000000000000010;
        16'b0000000110101101 : reciprocal = 16'b0000000000000010;
        16'b0000000110101110 : reciprocal = 16'b0000000000000010;
        16'b0000000110101111 : reciprocal = 16'b0000000000000010;
        16'b0000000110110000 : reciprocal = 16'b0000000000000010;
        16'b0000000110110001 : reciprocal = 16'b0000000000000010;
        16'b0000000110110010 : reciprocal = 16'b0000000000000010;
        16'b0000000110110011 : reciprocal = 16'b0000000000000010;
        16'b0000000110110100 : reciprocal = 16'b0000000000000010;
        16'b0000000110110101 : reciprocal = 16'b0000000000000010;
        16'b0000000110110110 : reciprocal = 16'b0000000000000010;
        16'b0000000110110111 : reciprocal = 16'b0000000000000010;
        16'b0000000110111000 : reciprocal = 16'b0000000000000010;
        16'b0000000110111001 : reciprocal = 16'b0000000000000010;
        16'b0000000110111010 : reciprocal = 16'b0000000000000010;
        16'b0000000110111011 : reciprocal = 16'b0000000000000010;
        16'b0000000110111100 : reciprocal = 16'b0000000000000010;
        16'b0000000110111101 : reciprocal = 16'b0000000000000010;
        16'b0000000110111110 : reciprocal = 16'b0000000000000010;
        16'b0000000110111111 : reciprocal = 16'b0000000000000010;
        16'b0000000111000000 : reciprocal = 16'b0000000000000010;
        16'b0000000111000001 : reciprocal = 16'b0000000000000010;
        16'b0000000111000010 : reciprocal = 16'b0000000000000010;
        16'b0000000111000011 : reciprocal = 16'b0000000000000010;
        16'b0000000111000100 : reciprocal = 16'b0000000000000010;
        16'b0000000111000101 : reciprocal = 16'b0000000000000010;
        16'b0000000111000110 : reciprocal = 16'b0000000000000010;
        16'b0000000111000111 : reciprocal = 16'b0000000000000010;
        16'b0000000111001000 : reciprocal = 16'b0000000000000010;
        16'b0000000111001001 : reciprocal = 16'b0000000000000010;
        16'b0000000111001010 : reciprocal = 16'b0000000000000010;
        16'b0000000111001011 : reciprocal = 16'b0000000000000010;
        16'b0000000111001100 : reciprocal = 16'b0000000000000010;
        16'b0000000111001101 : reciprocal = 16'b0000000000000010;
        16'b0000000111001110 : reciprocal = 16'b0000000000000010;
        16'b0000000111001111 : reciprocal = 16'b0000000000000010;
        16'b0000000111010000 : reciprocal = 16'b0000000000000010;
        16'b0000000111010001 : reciprocal = 16'b0000000000000010;
        16'b0000000111010010 : reciprocal = 16'b0000000000000010;
        16'b0000000111010011 : reciprocal = 16'b0000000000000010;
        16'b0000000111010100 : reciprocal = 16'b0000000000000010;
        16'b0000000111010101 : reciprocal = 16'b0000000000000010;
        16'b0000000111010110 : reciprocal = 16'b0000000000000010;
        16'b0000000111010111 : reciprocal = 16'b0000000000000010;
        16'b0000000111011000 : reciprocal = 16'b0000000000000010;
        16'b0000000111011001 : reciprocal = 16'b0000000000000010;
        16'b0000000111011010 : reciprocal = 16'b0000000000000010;
        16'b0000000111011011 : reciprocal = 16'b0000000000000010;
        16'b0000000111011100 : reciprocal = 16'b0000000000000010;
        16'b0000000111011101 : reciprocal = 16'b0000000000000010;
        16'b0000000111011110 : reciprocal = 16'b0000000000000010;
        16'b0000000111011111 : reciprocal = 16'b0000000000000010;
        16'b0000000111100000 : reciprocal = 16'b0000000000000010;
        16'b0000000111100001 : reciprocal = 16'b0000000000000010;
        16'b0000000111100010 : reciprocal = 16'b0000000000000010;
        16'b0000000111100011 : reciprocal = 16'b0000000000000010;
        16'b0000000111100100 : reciprocal = 16'b0000000000000010;
        16'b0000000111100101 : reciprocal = 16'b0000000000000010;
        16'b0000000111100110 : reciprocal = 16'b0000000000000010;
        16'b0000000111100111 : reciprocal = 16'b0000000000000010;
        16'b0000000111101000 : reciprocal = 16'b0000000000000010;
        16'b0000000111101001 : reciprocal = 16'b0000000000000010;
        16'b0000000111101010 : reciprocal = 16'b0000000000000010;
        16'b0000000111101011 : reciprocal = 16'b0000000000000010;
        16'b0000000111101100 : reciprocal = 16'b0000000000000010;
        16'b0000000111101101 : reciprocal = 16'b0000000000000010;
        16'b0000000111101110 : reciprocal = 16'b0000000000000010;
        16'b0000000111101111 : reciprocal = 16'b0000000000000010;
        16'b0000000111110000 : reciprocal = 16'b0000000000000010;
        16'b0000000111110001 : reciprocal = 16'b0000000000000010;
        16'b0000000111110010 : reciprocal = 16'b0000000000000010;
        16'b0000000111110011 : reciprocal = 16'b0000000000000010;
        16'b0000000111110100 : reciprocal = 16'b0000000000000010;
        16'b0000000111110101 : reciprocal = 16'b0000000000000010;
        16'b0000000111110110 : reciprocal = 16'b0000000000000010;
        16'b0000000111110111 : reciprocal = 16'b0000000000000010;
        16'b0000000111111000 : reciprocal = 16'b0000000000000010;
        16'b0000000111111001 : reciprocal = 16'b0000000000000010;
        16'b0000000111111010 : reciprocal = 16'b0000000000000010;
        16'b0000000111111011 : reciprocal = 16'b0000000000000010;
        16'b0000000111111100 : reciprocal = 16'b0000000000000010;
        16'b0000000111111101 : reciprocal = 16'b0000000000000010;
        16'b0000000111111110 : reciprocal = 16'b0000000000000010;
        16'b0000000111111111 : reciprocal = 16'b0000000000000010;
        16'b0000001000000000 : reciprocal = 16'b0000000000000010;
        16'b0000001000000001 : reciprocal = 16'b0000000000000010;
        16'b0000001000000010 : reciprocal = 16'b0000000000000010;
        16'b0000001000000011 : reciprocal = 16'b0000000000000010;
        16'b0000001000000100 : reciprocal = 16'b0000000000000010;
        16'b0000001000000101 : reciprocal = 16'b0000000000000010;
        16'b0000001000000110 : reciprocal = 16'b0000000000000010;
        16'b0000001000000111 : reciprocal = 16'b0000000000000010;
        16'b0000001000001000 : reciprocal = 16'b0000000000000010;
        16'b0000001000001001 : reciprocal = 16'b0000000000000010;
        16'b0000001000001010 : reciprocal = 16'b0000000000000010;
        16'b0000001000001011 : reciprocal = 16'b0000000000000010;
        16'b0000001000001100 : reciprocal = 16'b0000000000000010;
        16'b0000001000001101 : reciprocal = 16'b0000000000000010;
        16'b0000001000001110 : reciprocal = 16'b0000000000000010;
        16'b0000001000001111 : reciprocal = 16'b0000000000000010;
        16'b0000001000010000 : reciprocal = 16'b0000000000000010;
        16'b0000001000010001 : reciprocal = 16'b0000000000000010;
        16'b0000001000010010 : reciprocal = 16'b0000000000000010;
        16'b0000001000010011 : reciprocal = 16'b0000000000000010;
        16'b0000001000010100 : reciprocal = 16'b0000000000000010;
        16'b0000001000010101 : reciprocal = 16'b0000000000000010;
        16'b0000001000010110 : reciprocal = 16'b0000000000000010;
        16'b0000001000010111 : reciprocal = 16'b0000000000000010;
        16'b0000001000011000 : reciprocal = 16'b0000000000000010;
        16'b0000001000011001 : reciprocal = 16'b0000000000000010;
        16'b0000001000011010 : reciprocal = 16'b0000000000000010;
        16'b0000001000011011 : reciprocal = 16'b0000000000000010;
        16'b0000001000011100 : reciprocal = 16'b0000000000000010;
        16'b0000001000011101 : reciprocal = 16'b0000000000000010;
        16'b0000001000011110 : reciprocal = 16'b0000000000000010;
        16'b0000001000011111 : reciprocal = 16'b0000000000000010;
        16'b0000001000100000 : reciprocal = 16'b0000000000000010;
        16'b0000001000100001 : reciprocal = 16'b0000000000000010;
        16'b0000001000100010 : reciprocal = 16'b0000000000000010;
        16'b0000001000100011 : reciprocal = 16'b0000000000000010;
        16'b0000001000100100 : reciprocal = 16'b0000000000000010;
        16'b0000001000100101 : reciprocal = 16'b0000000000000010;
        16'b0000001000100110 : reciprocal = 16'b0000000000000010;
        16'b0000001000100111 : reciprocal = 16'b0000000000000010;
        16'b0000001000101000 : reciprocal = 16'b0000000000000010;
        16'b0000001000101001 : reciprocal = 16'b0000000000000010;
        16'b0000001000101010 : reciprocal = 16'b0000000000000010;
        16'b0000001000101011 : reciprocal = 16'b0000000000000010;
        16'b0000001000101100 : reciprocal = 16'b0000000000000010;
        16'b0000001000101101 : reciprocal = 16'b0000000000000010;
        16'b0000001000101110 : reciprocal = 16'b0000000000000010;
        16'b0000001000101111 : reciprocal = 16'b0000000000000010;
        16'b0000001000110000 : reciprocal = 16'b0000000000000010;
        16'b0000001000110001 : reciprocal = 16'b0000000000000010;
        16'b0000001000110010 : reciprocal = 16'b0000000000000010;
        16'b0000001000110011 : reciprocal = 16'b0000000000000010;
        16'b0000001000110100 : reciprocal = 16'b0000000000000010;
        16'b0000001000110101 : reciprocal = 16'b0000000000000010;
        16'b0000001000110110 : reciprocal = 16'b0000000000000010;
        16'b0000001000110111 : reciprocal = 16'b0000000000000010;
        16'b0000001000111000 : reciprocal = 16'b0000000000000010;
        16'b0000001000111001 : reciprocal = 16'b0000000000000010;
        16'b0000001000111010 : reciprocal = 16'b0000000000000010;
        16'b0000001000111011 : reciprocal = 16'b0000000000000010;
        16'b0000001000111100 : reciprocal = 16'b0000000000000010;
        16'b0000001000111101 : reciprocal = 16'b0000000000000010;
        16'b0000001000111110 : reciprocal = 16'b0000000000000010;
        16'b0000001000111111 : reciprocal = 16'b0000000000000010;
        16'b0000001001000000 : reciprocal = 16'b0000000000000010;
        16'b0000001001000001 : reciprocal = 16'b0000000000000010;
        16'b0000001001000010 : reciprocal = 16'b0000000000000010;
        16'b0000001001000011 : reciprocal = 16'b0000000000000010;
        16'b0000001001000100 : reciprocal = 16'b0000000000000010;
        16'b0000001001000101 : reciprocal = 16'b0000000000000010;
        16'b0000001001000110 : reciprocal = 16'b0000000000000010;
        16'b0000001001000111 : reciprocal = 16'b0000000000000010;
        16'b0000001001001000 : reciprocal = 16'b0000000000000010;
        16'b0000001001001001 : reciprocal = 16'b0000000000000010;
        16'b0000001001001010 : reciprocal = 16'b0000000000000010;
        16'b0000001001001011 : reciprocal = 16'b0000000000000010;
        16'b0000001001001100 : reciprocal = 16'b0000000000000010;
        16'b0000001001001101 : reciprocal = 16'b0000000000000010;
        16'b0000001001001110 : reciprocal = 16'b0000000000000010;
        16'b0000001001001111 : reciprocal = 16'b0000000000000010;
        16'b0000001001010000 : reciprocal = 16'b0000000000000010;
        16'b0000001001010001 : reciprocal = 16'b0000000000000010;
        16'b0000001001010010 : reciprocal = 16'b0000000000000010;
        16'b0000001001010011 : reciprocal = 16'b0000000000000010;
        16'b0000001001010100 : reciprocal = 16'b0000000000000010;
        16'b0000001001010101 : reciprocal = 16'b0000000000000010;
        16'b0000001001010110 : reciprocal = 16'b0000000000000010;
        16'b0000001001010111 : reciprocal = 16'b0000000000000010;
        16'b0000001001011000 : reciprocal = 16'b0000000000000010;
        16'b0000001001011001 : reciprocal = 16'b0000000000000010;
        16'b0000001001011010 : reciprocal = 16'b0000000000000010;
        16'b0000001001011011 : reciprocal = 16'b0000000000000010;
        16'b0000001001011100 : reciprocal = 16'b0000000000000010;
        16'b0000001001011101 : reciprocal = 16'b0000000000000010;
        16'b0000001001011110 : reciprocal = 16'b0000000000000010;
        16'b0000001001011111 : reciprocal = 16'b0000000000000010;
        16'b0000001001100000 : reciprocal = 16'b0000000000000010;
        16'b0000001001100001 : reciprocal = 16'b0000000000000010;
        16'b0000001001100010 : reciprocal = 16'b0000000000000010;
        16'b0000001001100011 : reciprocal = 16'b0000000000000010;
        16'b0000001001100100 : reciprocal = 16'b0000000000000010;
        16'b0000001001100101 : reciprocal = 16'b0000000000000010;
        16'b0000001001100110 : reciprocal = 16'b0000000000000010;
        16'b0000001001100111 : reciprocal = 16'b0000000000000010;
        16'b0000001001101000 : reciprocal = 16'b0000000000000010;
        16'b0000001001101001 : reciprocal = 16'b0000000000000010;
        16'b0000001001101010 : reciprocal = 16'b0000000000000010;
        16'b0000001001101011 : reciprocal = 16'b0000000000000010;
        16'b0000001001101100 : reciprocal = 16'b0000000000000010;
        16'b0000001001101101 : reciprocal = 16'b0000000000000010;
        16'b0000001001101110 : reciprocal = 16'b0000000000000010;
        16'b0000001001101111 : reciprocal = 16'b0000000000000010;
        16'b0000001001110000 : reciprocal = 16'b0000000000000010;
        16'b0000001001110001 : reciprocal = 16'b0000000000000010;
        16'b0000001001110010 : reciprocal = 16'b0000000000000010;
        16'b0000001001110011 : reciprocal = 16'b0000000000000010;
        16'b0000001001110100 : reciprocal = 16'b0000000000000010;
        16'b0000001001110101 : reciprocal = 16'b0000000000000010;
        16'b0000001001110110 : reciprocal = 16'b0000000000000010;
        16'b0000001001110111 : reciprocal = 16'b0000000000000010;
        16'b0000001001111000 : reciprocal = 16'b0000000000000010;
        16'b0000001001111001 : reciprocal = 16'b0000000000000010;
        16'b0000001001111010 : reciprocal = 16'b0000000000000010;
        16'b0000001001111011 : reciprocal = 16'b0000000000000010;
        16'b0000001001111100 : reciprocal = 16'b0000000000000010;
        16'b0000001001111101 : reciprocal = 16'b0000000000000010;
        16'b0000001001111110 : reciprocal = 16'b0000000000000010;
        16'b0000001001111111 : reciprocal = 16'b0000000000000010;
        16'b0000001010000000 : reciprocal = 16'b0000000000000010;
        16'b0000001010000001 : reciprocal = 16'b0000000000000010;
        16'b0000001010000010 : reciprocal = 16'b0000000000000010;
        16'b0000001010000011 : reciprocal = 16'b0000000000000010;
        16'b0000001010000100 : reciprocal = 16'b0000000000000010;
        16'b0000001010000101 : reciprocal = 16'b0000000000000010;
        16'b0000001010000110 : reciprocal = 16'b0000000000000010;
        16'b0000001010000111 : reciprocal = 16'b0000000000000010;
        16'b0000001010001000 : reciprocal = 16'b0000000000000010;
        16'b0000001010001001 : reciprocal = 16'b0000000000000010;
        16'b0000001010001010 : reciprocal = 16'b0000000000000010;
        16'b0000001010001011 : reciprocal = 16'b0000000000000010;
        16'b0000001010001100 : reciprocal = 16'b0000000000000010;
        16'b0000001010001101 : reciprocal = 16'b0000000000000010;
        16'b0000001010001110 : reciprocal = 16'b0000000000000010;
        16'b0000001010001111 : reciprocal = 16'b0000000000000010;
        16'b0000001010010000 : reciprocal = 16'b0000000000000010;
        16'b0000001010010001 : reciprocal = 16'b0000000000000010;
        16'b0000001010010010 : reciprocal = 16'b0000000000000010;
        16'b0000001010010011 : reciprocal = 16'b0000000000000010;
        16'b0000001010010100 : reciprocal = 16'b0000000000000010;
        16'b0000001010010101 : reciprocal = 16'b0000000000000010;
        16'b0000001010010110 : reciprocal = 16'b0000000000000010;
        16'b0000001010010111 : reciprocal = 16'b0000000000000010;
        16'b0000001010011000 : reciprocal = 16'b0000000000000010;
        16'b0000001010011001 : reciprocal = 16'b0000000000000010;
        16'b0000001010011010 : reciprocal = 16'b0000000000000010;
        16'b0000001010011011 : reciprocal = 16'b0000000000000010;
        16'b0000001010011100 : reciprocal = 16'b0000000000000010;
        16'b0000001010011101 : reciprocal = 16'b0000000000000010;
        16'b0000001010011110 : reciprocal = 16'b0000000000000010;
        16'b0000001010011111 : reciprocal = 16'b0000000000000010;
        16'b0000001010100000 : reciprocal = 16'b0000000000000010;
        16'b0000001010100001 : reciprocal = 16'b0000000000000010;
        16'b0000001010100010 : reciprocal = 16'b0000000000000010;
        16'b0000001010100011 : reciprocal = 16'b0000000000000010;
        16'b0000001010100100 : reciprocal = 16'b0000000000000010;
        16'b0000001010100101 : reciprocal = 16'b0000000000000010;
        16'b0000001010100110 : reciprocal = 16'b0000000000000010;
        16'b0000001010100111 : reciprocal = 16'b0000000000000010;
        16'b0000001010101000 : reciprocal = 16'b0000000000000010;
        16'b0000001010101001 : reciprocal = 16'b0000000000000010;
        16'b0000001010101010 : reciprocal = 16'b0000000000000010;
        16'b0000001010101011 : reciprocal = 16'b0000000000000001;
        16'b0000001010101100 : reciprocal = 16'b0000000000000001;
        16'b0000001010101101 : reciprocal = 16'b0000000000000001;
        16'b0000001010101110 : reciprocal = 16'b0000000000000001;
        16'b0000001010101111 : reciprocal = 16'b0000000000000001;
        16'b0000001010110000 : reciprocal = 16'b0000000000000001;
        16'b0000001010110001 : reciprocal = 16'b0000000000000001;
        16'b0000001010110010 : reciprocal = 16'b0000000000000001;
        16'b0000001010110011 : reciprocal = 16'b0000000000000001;
        16'b0000001010110100 : reciprocal = 16'b0000000000000001;
        16'b0000001010110101 : reciprocal = 16'b0000000000000001;
        16'b0000001010110110 : reciprocal = 16'b0000000000000001;
        16'b0000001010110111 : reciprocal = 16'b0000000000000001;
        16'b0000001010111000 : reciprocal = 16'b0000000000000001;
        16'b0000001010111001 : reciprocal = 16'b0000000000000001;
        16'b0000001010111010 : reciprocal = 16'b0000000000000001;
        16'b0000001010111011 : reciprocal = 16'b0000000000000001;
        16'b0000001010111100 : reciprocal = 16'b0000000000000001;
        16'b0000001010111101 : reciprocal = 16'b0000000000000001;
        16'b0000001010111110 : reciprocal = 16'b0000000000000001;
        16'b0000001010111111 : reciprocal = 16'b0000000000000001;
        16'b0000001011000000 : reciprocal = 16'b0000000000000001;
        16'b0000001011000001 : reciprocal = 16'b0000000000000001;
        16'b0000001011000010 : reciprocal = 16'b0000000000000001;
        16'b0000001011000011 : reciprocal = 16'b0000000000000001;
        16'b0000001011000100 : reciprocal = 16'b0000000000000001;
        16'b0000001011000101 : reciprocal = 16'b0000000000000001;
        16'b0000001011000110 : reciprocal = 16'b0000000000000001;
        16'b0000001011000111 : reciprocal = 16'b0000000000000001;
        16'b0000001011001000 : reciprocal = 16'b0000000000000001;
        16'b0000001011001001 : reciprocal = 16'b0000000000000001;
        16'b0000001011001010 : reciprocal = 16'b0000000000000001;
        16'b0000001011001011 : reciprocal = 16'b0000000000000001;
        16'b0000001011001100 : reciprocal = 16'b0000000000000001;
        16'b0000001011001101 : reciprocal = 16'b0000000000000001;
        16'b0000001011001110 : reciprocal = 16'b0000000000000001;
        16'b0000001011001111 : reciprocal = 16'b0000000000000001;
        16'b0000001011010000 : reciprocal = 16'b0000000000000001;
        16'b0000001011010001 : reciprocal = 16'b0000000000000001;
        16'b0000001011010010 : reciprocal = 16'b0000000000000001;
        16'b0000001011010011 : reciprocal = 16'b0000000000000001;
        16'b0000001011010100 : reciprocal = 16'b0000000000000001;
        16'b0000001011010101 : reciprocal = 16'b0000000000000001;
        16'b0000001011010110 : reciprocal = 16'b0000000000000001;
        16'b0000001011010111 : reciprocal = 16'b0000000000000001;
        16'b0000001011011000 : reciprocal = 16'b0000000000000001;
        16'b0000001011011001 : reciprocal = 16'b0000000000000001;
        16'b0000001011011010 : reciprocal = 16'b0000000000000001;
        16'b0000001011011011 : reciprocal = 16'b0000000000000001;
        16'b0000001011011100 : reciprocal = 16'b0000000000000001;
        16'b0000001011011101 : reciprocal = 16'b0000000000000001;
        16'b0000001011011110 : reciprocal = 16'b0000000000000001;
        16'b0000001011011111 : reciprocal = 16'b0000000000000001;
        16'b0000001011100000 : reciprocal = 16'b0000000000000001;
        16'b0000001011100001 : reciprocal = 16'b0000000000000001;
        16'b0000001011100010 : reciprocal = 16'b0000000000000001;
        16'b0000001011100011 : reciprocal = 16'b0000000000000001;
        16'b0000001011100100 : reciprocal = 16'b0000000000000001;
        16'b0000001011100101 : reciprocal = 16'b0000000000000001;
        16'b0000001011100110 : reciprocal = 16'b0000000000000001;
        16'b0000001011100111 : reciprocal = 16'b0000000000000001;
        16'b0000001011101000 : reciprocal = 16'b0000000000000001;
        16'b0000001011101001 : reciprocal = 16'b0000000000000001;
        16'b0000001011101010 : reciprocal = 16'b0000000000000001;
        16'b0000001011101011 : reciprocal = 16'b0000000000000001;
        16'b0000001011101100 : reciprocal = 16'b0000000000000001;
        16'b0000001011101101 : reciprocal = 16'b0000000000000001;
        16'b0000001011101110 : reciprocal = 16'b0000000000000001;
        16'b0000001011101111 : reciprocal = 16'b0000000000000001;
        16'b0000001011110000 : reciprocal = 16'b0000000000000001;
        16'b0000001011110001 : reciprocal = 16'b0000000000000001;
        16'b0000001011110010 : reciprocal = 16'b0000000000000001;
        16'b0000001011110011 : reciprocal = 16'b0000000000000001;
        16'b0000001011110100 : reciprocal = 16'b0000000000000001;
        16'b0000001011110101 : reciprocal = 16'b0000000000000001;
        16'b0000001011110110 : reciprocal = 16'b0000000000000001;
        16'b0000001011110111 : reciprocal = 16'b0000000000000001;
        16'b0000001011111000 : reciprocal = 16'b0000000000000001;
        16'b0000001011111001 : reciprocal = 16'b0000000000000001;
        16'b0000001011111010 : reciprocal = 16'b0000000000000001;
        16'b0000001011111011 : reciprocal = 16'b0000000000000001;
        16'b0000001011111100 : reciprocal = 16'b0000000000000001;
        16'b0000001011111101 : reciprocal = 16'b0000000000000001;
        16'b0000001011111110 : reciprocal = 16'b0000000000000001;
        16'b0000001011111111 : reciprocal = 16'b0000000000000001;
        16'b0000001100000000 : reciprocal = 16'b0000000000000001;
        16'b0000001100000001 : reciprocal = 16'b0000000000000001;
        16'b0000001100000010 : reciprocal = 16'b0000000000000001;
        16'b0000001100000011 : reciprocal = 16'b0000000000000001;
        16'b0000001100000100 : reciprocal = 16'b0000000000000001;
        16'b0000001100000101 : reciprocal = 16'b0000000000000001;
        16'b0000001100000110 : reciprocal = 16'b0000000000000001;
        16'b0000001100000111 : reciprocal = 16'b0000000000000001;
        16'b0000001100001000 : reciprocal = 16'b0000000000000001;
        16'b0000001100001001 : reciprocal = 16'b0000000000000001;
        16'b0000001100001010 : reciprocal = 16'b0000000000000001;
        16'b0000001100001011 : reciprocal = 16'b0000000000000001;
        16'b0000001100001100 : reciprocal = 16'b0000000000000001;
        16'b0000001100001101 : reciprocal = 16'b0000000000000001;
        16'b0000001100001110 : reciprocal = 16'b0000000000000001;
        16'b0000001100001111 : reciprocal = 16'b0000000000000001;
        16'b0000001100010000 : reciprocal = 16'b0000000000000001;
        16'b0000001100010001 : reciprocal = 16'b0000000000000001;
        16'b0000001100010010 : reciprocal = 16'b0000000000000001;
        16'b0000001100010011 : reciprocal = 16'b0000000000000001;
        16'b0000001100010100 : reciprocal = 16'b0000000000000001;
        16'b0000001100010101 : reciprocal = 16'b0000000000000001;
        16'b0000001100010110 : reciprocal = 16'b0000000000000001;
        16'b0000001100010111 : reciprocal = 16'b0000000000000001;
        16'b0000001100011000 : reciprocal = 16'b0000000000000001;
        16'b0000001100011001 : reciprocal = 16'b0000000000000001;
        16'b0000001100011010 : reciprocal = 16'b0000000000000001;
        16'b0000001100011011 : reciprocal = 16'b0000000000000001;
        16'b0000001100011100 : reciprocal = 16'b0000000000000001;
        16'b0000001100011101 : reciprocal = 16'b0000000000000001;
        16'b0000001100011110 : reciprocal = 16'b0000000000000001;
        16'b0000001100011111 : reciprocal = 16'b0000000000000001;
        16'b0000001100100000 : reciprocal = 16'b0000000000000001;
        16'b0000001100100001 : reciprocal = 16'b0000000000000001;
        16'b0000001100100010 : reciprocal = 16'b0000000000000001;
        16'b0000001100100011 : reciprocal = 16'b0000000000000001;
        16'b0000001100100100 : reciprocal = 16'b0000000000000001;
        16'b0000001100100101 : reciprocal = 16'b0000000000000001;
        16'b0000001100100110 : reciprocal = 16'b0000000000000001;
        16'b0000001100100111 : reciprocal = 16'b0000000000000001;
        16'b0000001100101000 : reciprocal = 16'b0000000000000001;
        16'b0000001100101001 : reciprocal = 16'b0000000000000001;
        16'b0000001100101010 : reciprocal = 16'b0000000000000001;
        16'b0000001100101011 : reciprocal = 16'b0000000000000001;
        16'b0000001100101100 : reciprocal = 16'b0000000000000001;
        16'b0000001100101101 : reciprocal = 16'b0000000000000001;
        16'b0000001100101110 : reciprocal = 16'b0000000000000001;
        16'b0000001100101111 : reciprocal = 16'b0000000000000001;
        16'b0000001100110000 : reciprocal = 16'b0000000000000001;
        16'b0000001100110001 : reciprocal = 16'b0000000000000001;
        16'b0000001100110010 : reciprocal = 16'b0000000000000001;
        16'b0000001100110011 : reciprocal = 16'b0000000000000001;
        16'b0000001100110100 : reciprocal = 16'b0000000000000001;
        16'b0000001100110101 : reciprocal = 16'b0000000000000001;
        16'b0000001100110110 : reciprocal = 16'b0000000000000001;
        16'b0000001100110111 : reciprocal = 16'b0000000000000001;
        16'b0000001100111000 : reciprocal = 16'b0000000000000001;
        16'b0000001100111001 : reciprocal = 16'b0000000000000001;
        16'b0000001100111010 : reciprocal = 16'b0000000000000001;
        16'b0000001100111011 : reciprocal = 16'b0000000000000001;
        16'b0000001100111100 : reciprocal = 16'b0000000000000001;
        16'b0000001100111101 : reciprocal = 16'b0000000000000001;
        16'b0000001100111110 : reciprocal = 16'b0000000000000001;
        16'b0000001100111111 : reciprocal = 16'b0000000000000001;
        16'b0000001101000000 : reciprocal = 16'b0000000000000001;
        16'b0000001101000001 : reciprocal = 16'b0000000000000001;
        16'b0000001101000010 : reciprocal = 16'b0000000000000001;
        16'b0000001101000011 : reciprocal = 16'b0000000000000001;
        16'b0000001101000100 : reciprocal = 16'b0000000000000001;
        16'b0000001101000101 : reciprocal = 16'b0000000000000001;
        16'b0000001101000110 : reciprocal = 16'b0000000000000001;
        16'b0000001101000111 : reciprocal = 16'b0000000000000001;
        16'b0000001101001000 : reciprocal = 16'b0000000000000001;
        16'b0000001101001001 : reciprocal = 16'b0000000000000001;
        16'b0000001101001010 : reciprocal = 16'b0000000000000001;
        16'b0000001101001011 : reciprocal = 16'b0000000000000001;
        16'b0000001101001100 : reciprocal = 16'b0000000000000001;
        16'b0000001101001101 : reciprocal = 16'b0000000000000001;
        16'b0000001101001110 : reciprocal = 16'b0000000000000001;
        16'b0000001101001111 : reciprocal = 16'b0000000000000001;
        16'b0000001101010000 : reciprocal = 16'b0000000000000001;
        16'b0000001101010001 : reciprocal = 16'b0000000000000001;
        16'b0000001101010010 : reciprocal = 16'b0000000000000001;
        16'b0000001101010011 : reciprocal = 16'b0000000000000001;
        16'b0000001101010100 : reciprocal = 16'b0000000000000001;
        16'b0000001101010101 : reciprocal = 16'b0000000000000001;
        16'b0000001101010110 : reciprocal = 16'b0000000000000001;
        16'b0000001101010111 : reciprocal = 16'b0000000000000001;
        16'b0000001101011000 : reciprocal = 16'b0000000000000001;
        16'b0000001101011001 : reciprocal = 16'b0000000000000001;
        16'b0000001101011010 : reciprocal = 16'b0000000000000001;
        16'b0000001101011011 : reciprocal = 16'b0000000000000001;
        16'b0000001101011100 : reciprocal = 16'b0000000000000001;
        16'b0000001101011101 : reciprocal = 16'b0000000000000001;
        16'b0000001101011110 : reciprocal = 16'b0000000000000001;
        16'b0000001101011111 : reciprocal = 16'b0000000000000001;
        16'b0000001101100000 : reciprocal = 16'b0000000000000001;
        16'b0000001101100001 : reciprocal = 16'b0000000000000001;
        16'b0000001101100010 : reciprocal = 16'b0000000000000001;
        16'b0000001101100011 : reciprocal = 16'b0000000000000001;
        16'b0000001101100100 : reciprocal = 16'b0000000000000001;
        16'b0000001101100101 : reciprocal = 16'b0000000000000001;
        16'b0000001101100110 : reciprocal = 16'b0000000000000001;
        16'b0000001101100111 : reciprocal = 16'b0000000000000001;
        16'b0000001101101000 : reciprocal = 16'b0000000000000001;
        16'b0000001101101001 : reciprocal = 16'b0000000000000001;
        16'b0000001101101010 : reciprocal = 16'b0000000000000001;
        16'b0000001101101011 : reciprocal = 16'b0000000000000001;
        16'b0000001101101100 : reciprocal = 16'b0000000000000001;
        16'b0000001101101101 : reciprocal = 16'b0000000000000001;
        16'b0000001101101110 : reciprocal = 16'b0000000000000001;
        16'b0000001101101111 : reciprocal = 16'b0000000000000001;
        16'b0000001101110000 : reciprocal = 16'b0000000000000001;
        16'b0000001101110001 : reciprocal = 16'b0000000000000001;
        16'b0000001101110010 : reciprocal = 16'b0000000000000001;
        16'b0000001101110011 : reciprocal = 16'b0000000000000001;
        16'b0000001101110100 : reciprocal = 16'b0000000000000001;
        16'b0000001101110101 : reciprocal = 16'b0000000000000001;
        16'b0000001101110110 : reciprocal = 16'b0000000000000001;
        16'b0000001101110111 : reciprocal = 16'b0000000000000001;
        16'b0000001101111000 : reciprocal = 16'b0000000000000001;
        16'b0000001101111001 : reciprocal = 16'b0000000000000001;
        16'b0000001101111010 : reciprocal = 16'b0000000000000001;
        16'b0000001101111011 : reciprocal = 16'b0000000000000001;
        16'b0000001101111100 : reciprocal = 16'b0000000000000001;
        16'b0000001101111101 : reciprocal = 16'b0000000000000001;
        16'b0000001101111110 : reciprocal = 16'b0000000000000001;
        16'b0000001101111111 : reciprocal = 16'b0000000000000001;
        16'b0000001110000000 : reciprocal = 16'b0000000000000001;
        16'b0000001110000001 : reciprocal = 16'b0000000000000001;
        16'b0000001110000010 : reciprocal = 16'b0000000000000001;
        16'b0000001110000011 : reciprocal = 16'b0000000000000001;
        16'b0000001110000100 : reciprocal = 16'b0000000000000001;
        16'b0000001110000101 : reciprocal = 16'b0000000000000001;
        16'b0000001110000110 : reciprocal = 16'b0000000000000001;
        16'b0000001110000111 : reciprocal = 16'b0000000000000001;
        16'b0000001110001000 : reciprocal = 16'b0000000000000001;
        16'b0000001110001001 : reciprocal = 16'b0000000000000001;
        16'b0000001110001010 : reciprocal = 16'b0000000000000001;
        16'b0000001110001011 : reciprocal = 16'b0000000000000001;
        16'b0000001110001100 : reciprocal = 16'b0000000000000001;
        16'b0000001110001101 : reciprocal = 16'b0000000000000001;
        16'b0000001110001110 : reciprocal = 16'b0000000000000001;
        16'b0000001110001111 : reciprocal = 16'b0000000000000001;
        16'b0000001110010000 : reciprocal = 16'b0000000000000001;
        16'b0000001110010001 : reciprocal = 16'b0000000000000001;
        16'b0000001110010010 : reciprocal = 16'b0000000000000001;
        16'b0000001110010011 : reciprocal = 16'b0000000000000001;
        16'b0000001110010100 : reciprocal = 16'b0000000000000001;
        16'b0000001110010101 : reciprocal = 16'b0000000000000001;
        16'b0000001110010110 : reciprocal = 16'b0000000000000001;
        16'b0000001110010111 : reciprocal = 16'b0000000000000001;
        16'b0000001110011000 : reciprocal = 16'b0000000000000001;
        16'b0000001110011001 : reciprocal = 16'b0000000000000001;
        16'b0000001110011010 : reciprocal = 16'b0000000000000001;
        16'b0000001110011011 : reciprocal = 16'b0000000000000001;
        16'b0000001110011100 : reciprocal = 16'b0000000000000001;
        16'b0000001110011101 : reciprocal = 16'b0000000000000001;
        16'b0000001110011110 : reciprocal = 16'b0000000000000001;
        16'b0000001110011111 : reciprocal = 16'b0000000000000001;
        16'b0000001110100000 : reciprocal = 16'b0000000000000001;
        16'b0000001110100001 : reciprocal = 16'b0000000000000001;
        16'b0000001110100010 : reciprocal = 16'b0000000000000001;
        16'b0000001110100011 : reciprocal = 16'b0000000000000001;
        16'b0000001110100100 : reciprocal = 16'b0000000000000001;
        16'b0000001110100101 : reciprocal = 16'b0000000000000001;
        16'b0000001110100110 : reciprocal = 16'b0000000000000001;
        16'b0000001110100111 : reciprocal = 16'b0000000000000001;
        16'b0000001110101000 : reciprocal = 16'b0000000000000001;
        16'b0000001110101001 : reciprocal = 16'b0000000000000001;
        16'b0000001110101010 : reciprocal = 16'b0000000000000001;
        16'b0000001110101011 : reciprocal = 16'b0000000000000001;
        16'b0000001110101100 : reciprocal = 16'b0000000000000001;
        16'b0000001110101101 : reciprocal = 16'b0000000000000001;
        16'b0000001110101110 : reciprocal = 16'b0000000000000001;
        16'b0000001110101111 : reciprocal = 16'b0000000000000001;
        16'b0000001110110000 : reciprocal = 16'b0000000000000001;
        16'b0000001110110001 : reciprocal = 16'b0000000000000001;
        16'b0000001110110010 : reciprocal = 16'b0000000000000001;
        16'b0000001110110011 : reciprocal = 16'b0000000000000001;
        16'b0000001110110100 : reciprocal = 16'b0000000000000001;
        16'b0000001110110101 : reciprocal = 16'b0000000000000001;
        16'b0000001110110110 : reciprocal = 16'b0000000000000001;
        16'b0000001110110111 : reciprocal = 16'b0000000000000001;
        16'b0000001110111000 : reciprocal = 16'b0000000000000001;
        16'b0000001110111001 : reciprocal = 16'b0000000000000001;
        16'b0000001110111010 : reciprocal = 16'b0000000000000001;
        16'b0000001110111011 : reciprocal = 16'b0000000000000001;
        16'b0000001110111100 : reciprocal = 16'b0000000000000001;
        16'b0000001110111101 : reciprocal = 16'b0000000000000001;
        16'b0000001110111110 : reciprocal = 16'b0000000000000001;
        16'b0000001110111111 : reciprocal = 16'b0000000000000001;
        16'b0000001111000000 : reciprocal = 16'b0000000000000001;
        16'b0000001111000001 : reciprocal = 16'b0000000000000001;
        16'b0000001111000010 : reciprocal = 16'b0000000000000001;
        16'b0000001111000011 : reciprocal = 16'b0000000000000001;
        16'b0000001111000100 : reciprocal = 16'b0000000000000001;
        16'b0000001111000101 : reciprocal = 16'b0000000000000001;
        16'b0000001111000110 : reciprocal = 16'b0000000000000001;
        16'b0000001111000111 : reciprocal = 16'b0000000000000001;
        16'b0000001111001000 : reciprocal = 16'b0000000000000001;
        16'b0000001111001001 : reciprocal = 16'b0000000000000001;
        16'b0000001111001010 : reciprocal = 16'b0000000000000001;
        16'b0000001111001011 : reciprocal = 16'b0000000000000001;
        16'b0000001111001100 : reciprocal = 16'b0000000000000001;
        16'b0000001111001101 : reciprocal = 16'b0000000000000001;
        16'b0000001111001110 : reciprocal = 16'b0000000000000001;
        16'b0000001111001111 : reciprocal = 16'b0000000000000001;
        16'b0000001111010000 : reciprocal = 16'b0000000000000001;
        16'b0000001111010001 : reciprocal = 16'b0000000000000001;
        16'b0000001111010010 : reciprocal = 16'b0000000000000001;
        16'b0000001111010011 : reciprocal = 16'b0000000000000001;
        16'b0000001111010100 : reciprocal = 16'b0000000000000001;
        16'b0000001111010101 : reciprocal = 16'b0000000000000001;
        16'b0000001111010110 : reciprocal = 16'b0000000000000001;
        16'b0000001111010111 : reciprocal = 16'b0000000000000001;
        16'b0000001111011000 : reciprocal = 16'b0000000000000001;
        16'b0000001111011001 : reciprocal = 16'b0000000000000001;
        16'b0000001111011010 : reciprocal = 16'b0000000000000001;
        16'b0000001111011011 : reciprocal = 16'b0000000000000001;
        16'b0000001111011100 : reciprocal = 16'b0000000000000001;
        16'b0000001111011101 : reciprocal = 16'b0000000000000001;
        16'b0000001111011110 : reciprocal = 16'b0000000000000001;
        16'b0000001111011111 : reciprocal = 16'b0000000000000001;
        16'b0000001111100000 : reciprocal = 16'b0000000000000001;
        16'b0000001111100001 : reciprocal = 16'b0000000000000001;
        16'b0000001111100010 : reciprocal = 16'b0000000000000001;
        16'b0000001111100011 : reciprocal = 16'b0000000000000001;
        16'b0000001111100100 : reciprocal = 16'b0000000000000001;
        16'b0000001111100101 : reciprocal = 16'b0000000000000001;
        16'b0000001111100110 : reciprocal = 16'b0000000000000001;
        16'b0000001111100111 : reciprocal = 16'b0000000000000001;
        16'b0000001111101000 : reciprocal = 16'b0000000000000001;
        16'b0000001111101001 : reciprocal = 16'b0000000000000001;
        16'b0000001111101010 : reciprocal = 16'b0000000000000001;
        16'b0000001111101011 : reciprocal = 16'b0000000000000001;
        16'b0000001111101100 : reciprocal = 16'b0000000000000001;
        16'b0000001111101101 : reciprocal = 16'b0000000000000001;
        16'b0000001111101110 : reciprocal = 16'b0000000000000001;
        16'b0000001111101111 : reciprocal = 16'b0000000000000001;
        16'b0000001111110000 : reciprocal = 16'b0000000000000001;
        16'b0000001111110001 : reciprocal = 16'b0000000000000001;
        16'b0000001111110010 : reciprocal = 16'b0000000000000001;
        16'b0000001111110011 : reciprocal = 16'b0000000000000001;
        16'b0000001111110100 : reciprocal = 16'b0000000000000001;
        16'b0000001111110101 : reciprocal = 16'b0000000000000001;
        16'b0000001111110110 : reciprocal = 16'b0000000000000001;
        16'b0000001111110111 : reciprocal = 16'b0000000000000001;
        16'b0000001111111000 : reciprocal = 16'b0000000000000001;
        16'b0000001111111001 : reciprocal = 16'b0000000000000001;
        16'b0000001111111010 : reciprocal = 16'b0000000000000001;
        16'b0000001111111011 : reciprocal = 16'b0000000000000001;
        16'b0000001111111100 : reciprocal = 16'b0000000000000001;
        16'b0000001111111101 : reciprocal = 16'b0000000000000001;
        16'b0000001111111110 : reciprocal = 16'b0000000000000001;
        16'b0000001111111111 : reciprocal = 16'b0000000000000001;
        16'b0000010000000000 : reciprocal = 16'b0000000000000001;
        16'b0000010000000001 : reciprocal = 16'b0000000000000001;
        16'b0000010000000010 : reciprocal = 16'b0000000000000001;
        16'b0000010000000011 : reciprocal = 16'b0000000000000001;
        16'b0000010000000100 : reciprocal = 16'b0000000000000001;
        16'b0000010000000101 : reciprocal = 16'b0000000000000001;
        16'b0000010000000110 : reciprocal = 16'b0000000000000001;
        16'b0000010000000111 : reciprocal = 16'b0000000000000001;
        16'b0000010000001000 : reciprocal = 16'b0000000000000001;
        16'b0000010000001001 : reciprocal = 16'b0000000000000001;
        16'b0000010000001010 : reciprocal = 16'b0000000000000001;
        16'b0000010000001011 : reciprocal = 16'b0000000000000001;
        16'b0000010000001100 : reciprocal = 16'b0000000000000001;
        16'b0000010000001101 : reciprocal = 16'b0000000000000001;
        16'b0000010000001110 : reciprocal = 16'b0000000000000001;
        16'b0000010000001111 : reciprocal = 16'b0000000000000001;
        16'b0000010000010000 : reciprocal = 16'b0000000000000001;
        16'b0000010000010001 : reciprocal = 16'b0000000000000001;
        16'b0000010000010010 : reciprocal = 16'b0000000000000001;
        16'b0000010000010011 : reciprocal = 16'b0000000000000001;
        16'b0000010000010100 : reciprocal = 16'b0000000000000001;
        16'b0000010000010101 : reciprocal = 16'b0000000000000001;
        16'b0000010000010110 : reciprocal = 16'b0000000000000001;
        16'b0000010000010111 : reciprocal = 16'b0000000000000001;
        16'b0000010000011000 : reciprocal = 16'b0000000000000001;
        16'b0000010000011001 : reciprocal = 16'b0000000000000001;
        16'b0000010000011010 : reciprocal = 16'b0000000000000001;
        16'b0000010000011011 : reciprocal = 16'b0000000000000001;
        16'b0000010000011100 : reciprocal = 16'b0000000000000001;
        16'b0000010000011101 : reciprocal = 16'b0000000000000001;
        16'b0000010000011110 : reciprocal = 16'b0000000000000001;
        16'b0000010000011111 : reciprocal = 16'b0000000000000001;
        16'b0000010000100000 : reciprocal = 16'b0000000000000001;
        16'b0000010000100001 : reciprocal = 16'b0000000000000001;
        16'b0000010000100010 : reciprocal = 16'b0000000000000001;
        16'b0000010000100011 : reciprocal = 16'b0000000000000001;
        16'b0000010000100100 : reciprocal = 16'b0000000000000001;
        16'b0000010000100101 : reciprocal = 16'b0000000000000001;
        16'b0000010000100110 : reciprocal = 16'b0000000000000001;
        16'b0000010000100111 : reciprocal = 16'b0000000000000001;
        16'b0000010000101000 : reciprocal = 16'b0000000000000001;
        16'b0000010000101001 : reciprocal = 16'b0000000000000001;
        16'b0000010000101010 : reciprocal = 16'b0000000000000001;
        16'b0000010000101011 : reciprocal = 16'b0000000000000001;
        16'b0000010000101100 : reciprocal = 16'b0000000000000001;
        16'b0000010000101101 : reciprocal = 16'b0000000000000001;
        16'b0000010000101110 : reciprocal = 16'b0000000000000001;
        16'b0000010000101111 : reciprocal = 16'b0000000000000001;
        16'b0000010000110000 : reciprocal = 16'b0000000000000001;
        16'b0000010000110001 : reciprocal = 16'b0000000000000001;
        16'b0000010000110010 : reciprocal = 16'b0000000000000001;
        16'b0000010000110011 : reciprocal = 16'b0000000000000001;
        16'b0000010000110100 : reciprocal = 16'b0000000000000001;
        16'b0000010000110101 : reciprocal = 16'b0000000000000001;
        16'b0000010000110110 : reciprocal = 16'b0000000000000001;
        16'b0000010000110111 : reciprocal = 16'b0000000000000001;
        16'b0000010000111000 : reciprocal = 16'b0000000000000001;
        16'b0000010000111001 : reciprocal = 16'b0000000000000001;
        16'b0000010000111010 : reciprocal = 16'b0000000000000001;
        16'b0000010000111011 : reciprocal = 16'b0000000000000001;
        16'b0000010000111100 : reciprocal = 16'b0000000000000001;
        16'b0000010000111101 : reciprocal = 16'b0000000000000001;
        16'b0000010000111110 : reciprocal = 16'b0000000000000001;
        16'b0000010000111111 : reciprocal = 16'b0000000000000001;
        16'b0000010001000000 : reciprocal = 16'b0000000000000001;
        16'b0000010001000001 : reciprocal = 16'b0000000000000001;
        16'b0000010001000010 : reciprocal = 16'b0000000000000001;
        16'b0000010001000011 : reciprocal = 16'b0000000000000001;
        16'b0000010001000100 : reciprocal = 16'b0000000000000001;
        16'b0000010001000101 : reciprocal = 16'b0000000000000001;
        16'b0000010001000110 : reciprocal = 16'b0000000000000001;
        16'b0000010001000111 : reciprocal = 16'b0000000000000001;
        16'b0000010001001000 : reciprocal = 16'b0000000000000001;
        16'b0000010001001001 : reciprocal = 16'b0000000000000001;
        16'b0000010001001010 : reciprocal = 16'b0000000000000001;
        16'b0000010001001011 : reciprocal = 16'b0000000000000001;
        16'b0000010001001100 : reciprocal = 16'b0000000000000001;
        16'b0000010001001101 : reciprocal = 16'b0000000000000001;
        16'b0000010001001110 : reciprocal = 16'b0000000000000001;
        16'b0000010001001111 : reciprocal = 16'b0000000000000001;
        16'b0000010001010000 : reciprocal = 16'b0000000000000001;
        16'b0000010001010001 : reciprocal = 16'b0000000000000001;
        16'b0000010001010010 : reciprocal = 16'b0000000000000001;
        16'b0000010001010011 : reciprocal = 16'b0000000000000001;
        16'b0000010001010100 : reciprocal = 16'b0000000000000001;
        16'b0000010001010101 : reciprocal = 16'b0000000000000001;
        16'b0000010001010110 : reciprocal = 16'b0000000000000001;
        16'b0000010001010111 : reciprocal = 16'b0000000000000001;
        16'b0000010001011000 : reciprocal = 16'b0000000000000001;
        16'b0000010001011001 : reciprocal = 16'b0000000000000001;
        16'b0000010001011010 : reciprocal = 16'b0000000000000001;
        16'b0000010001011011 : reciprocal = 16'b0000000000000001;
        16'b0000010001011100 : reciprocal = 16'b0000000000000001;
        16'b0000010001011101 : reciprocal = 16'b0000000000000001;
        16'b0000010001011110 : reciprocal = 16'b0000000000000001;
        16'b0000010001011111 : reciprocal = 16'b0000000000000001;
        16'b0000010001100000 : reciprocal = 16'b0000000000000001;
        16'b0000010001100001 : reciprocal = 16'b0000000000000001;
        16'b0000010001100010 : reciprocal = 16'b0000000000000001;
        16'b0000010001100011 : reciprocal = 16'b0000000000000001;
        16'b0000010001100100 : reciprocal = 16'b0000000000000001;
        16'b0000010001100101 : reciprocal = 16'b0000000000000001;
        16'b0000010001100110 : reciprocal = 16'b0000000000000001;
        16'b0000010001100111 : reciprocal = 16'b0000000000000001;
        16'b0000010001101000 : reciprocal = 16'b0000000000000001;
        16'b0000010001101001 : reciprocal = 16'b0000000000000001;
        16'b0000010001101010 : reciprocal = 16'b0000000000000001;
        16'b0000010001101011 : reciprocal = 16'b0000000000000001;
        16'b0000010001101100 : reciprocal = 16'b0000000000000001;
        16'b0000010001101101 : reciprocal = 16'b0000000000000001;
        16'b0000010001101110 : reciprocal = 16'b0000000000000001;
        16'b0000010001101111 : reciprocal = 16'b0000000000000001;
        16'b0000010001110000 : reciprocal = 16'b0000000000000001;
        16'b0000010001110001 : reciprocal = 16'b0000000000000001;
        16'b0000010001110010 : reciprocal = 16'b0000000000000001;
        16'b0000010001110011 : reciprocal = 16'b0000000000000001;
        16'b0000010001110100 : reciprocal = 16'b0000000000000001;
        16'b0000010001110101 : reciprocal = 16'b0000000000000001;
        16'b0000010001110110 : reciprocal = 16'b0000000000000001;
        16'b0000010001110111 : reciprocal = 16'b0000000000000001;
        16'b0000010001111000 : reciprocal = 16'b0000000000000001;
        16'b0000010001111001 : reciprocal = 16'b0000000000000001;
        16'b0000010001111010 : reciprocal = 16'b0000000000000001;
        16'b0000010001111011 : reciprocal = 16'b0000000000000001;
        16'b0000010001111100 : reciprocal = 16'b0000000000000001;
        16'b0000010001111101 : reciprocal = 16'b0000000000000001;
        16'b0000010001111110 : reciprocal = 16'b0000000000000001;
        16'b0000010001111111 : reciprocal = 16'b0000000000000001;
        16'b0000010010000000 : reciprocal = 16'b0000000000000001;
        16'b0000010010000001 : reciprocal = 16'b0000000000000001;
        16'b0000010010000010 : reciprocal = 16'b0000000000000001;
        16'b0000010010000011 : reciprocal = 16'b0000000000000001;
        16'b0000010010000100 : reciprocal = 16'b0000000000000001;
        16'b0000010010000101 : reciprocal = 16'b0000000000000001;
        16'b0000010010000110 : reciprocal = 16'b0000000000000001;
        16'b0000010010000111 : reciprocal = 16'b0000000000000001;
        16'b0000010010001000 : reciprocal = 16'b0000000000000001;
        16'b0000010010001001 : reciprocal = 16'b0000000000000001;
        16'b0000010010001010 : reciprocal = 16'b0000000000000001;
        16'b0000010010001011 : reciprocal = 16'b0000000000000001;
        16'b0000010010001100 : reciprocal = 16'b0000000000000001;
        16'b0000010010001101 : reciprocal = 16'b0000000000000001;
        16'b0000010010001110 : reciprocal = 16'b0000000000000001;
        16'b0000010010001111 : reciprocal = 16'b0000000000000001;
        16'b0000010010010000 : reciprocal = 16'b0000000000000001;
        16'b0000010010010001 : reciprocal = 16'b0000000000000001;
        16'b0000010010010010 : reciprocal = 16'b0000000000000001;
        16'b0000010010010011 : reciprocal = 16'b0000000000000001;
        16'b0000010010010100 : reciprocal = 16'b0000000000000001;
        16'b0000010010010101 : reciprocal = 16'b0000000000000001;
        16'b0000010010010110 : reciprocal = 16'b0000000000000001;
        16'b0000010010010111 : reciprocal = 16'b0000000000000001;
        16'b0000010010011000 : reciprocal = 16'b0000000000000001;
        16'b0000010010011001 : reciprocal = 16'b0000000000000001;
        16'b0000010010011010 : reciprocal = 16'b0000000000000001;
        16'b0000010010011011 : reciprocal = 16'b0000000000000001;
        16'b0000010010011100 : reciprocal = 16'b0000000000000001;
        16'b0000010010011101 : reciprocal = 16'b0000000000000001;
        16'b0000010010011110 : reciprocal = 16'b0000000000000001;
        16'b0000010010011111 : reciprocal = 16'b0000000000000001;
        16'b0000010010100000 : reciprocal = 16'b0000000000000001;
        16'b0000010010100001 : reciprocal = 16'b0000000000000001;
        16'b0000010010100010 : reciprocal = 16'b0000000000000001;
        16'b0000010010100011 : reciprocal = 16'b0000000000000001;
        16'b0000010010100100 : reciprocal = 16'b0000000000000001;
        16'b0000010010100101 : reciprocal = 16'b0000000000000001;
        16'b0000010010100110 : reciprocal = 16'b0000000000000001;
        16'b0000010010100111 : reciprocal = 16'b0000000000000001;
        16'b0000010010101000 : reciprocal = 16'b0000000000000001;
        16'b0000010010101001 : reciprocal = 16'b0000000000000001;
        16'b0000010010101010 : reciprocal = 16'b0000000000000001;
        16'b0000010010101011 : reciprocal = 16'b0000000000000001;
        16'b0000010010101100 : reciprocal = 16'b0000000000000001;
        16'b0000010010101101 : reciprocal = 16'b0000000000000001;
        16'b0000010010101110 : reciprocal = 16'b0000000000000001;
        16'b0000010010101111 : reciprocal = 16'b0000000000000001;
        16'b0000010010110000 : reciprocal = 16'b0000000000000001;
        16'b0000010010110001 : reciprocal = 16'b0000000000000001;
        16'b0000010010110010 : reciprocal = 16'b0000000000000001;
        16'b0000010010110011 : reciprocal = 16'b0000000000000001;
        16'b0000010010110100 : reciprocal = 16'b0000000000000001;
        16'b0000010010110101 : reciprocal = 16'b0000000000000001;
        16'b0000010010110110 : reciprocal = 16'b0000000000000001;
        16'b0000010010110111 : reciprocal = 16'b0000000000000001;
        16'b0000010010111000 : reciprocal = 16'b0000000000000001;
        16'b0000010010111001 : reciprocal = 16'b0000000000000001;
        16'b0000010010111010 : reciprocal = 16'b0000000000000001;
        16'b0000010010111011 : reciprocal = 16'b0000000000000001;
        16'b0000010010111100 : reciprocal = 16'b0000000000000001;
        16'b0000010010111101 : reciprocal = 16'b0000000000000001;
        16'b0000010010111110 : reciprocal = 16'b0000000000000001;
        16'b0000010010111111 : reciprocal = 16'b0000000000000001;
        16'b0000010011000000 : reciprocal = 16'b0000000000000001;
        16'b0000010011000001 : reciprocal = 16'b0000000000000001;
        16'b0000010011000010 : reciprocal = 16'b0000000000000001;
        16'b0000010011000011 : reciprocal = 16'b0000000000000001;
        16'b0000010011000100 : reciprocal = 16'b0000000000000001;
        16'b0000010011000101 : reciprocal = 16'b0000000000000001;
        16'b0000010011000110 : reciprocal = 16'b0000000000000001;
        16'b0000010011000111 : reciprocal = 16'b0000000000000001;
        16'b0000010011001000 : reciprocal = 16'b0000000000000001;
        16'b0000010011001001 : reciprocal = 16'b0000000000000001;
        16'b0000010011001010 : reciprocal = 16'b0000000000000001;
        16'b0000010011001011 : reciprocal = 16'b0000000000000001;
        16'b0000010011001100 : reciprocal = 16'b0000000000000001;
        16'b0000010011001101 : reciprocal = 16'b0000000000000001;
        16'b0000010011001110 : reciprocal = 16'b0000000000000001;
        16'b0000010011001111 : reciprocal = 16'b0000000000000001;
        16'b0000010011010000 : reciprocal = 16'b0000000000000001;
        16'b0000010011010001 : reciprocal = 16'b0000000000000001;
        16'b0000010011010010 : reciprocal = 16'b0000000000000001;
        16'b0000010011010011 : reciprocal = 16'b0000000000000001;
        16'b0000010011010100 : reciprocal = 16'b0000000000000001;
        16'b0000010011010101 : reciprocal = 16'b0000000000000001;
        16'b0000010011010110 : reciprocal = 16'b0000000000000001;
        16'b0000010011010111 : reciprocal = 16'b0000000000000001;
        16'b0000010011011000 : reciprocal = 16'b0000000000000001;
        16'b0000010011011001 : reciprocal = 16'b0000000000000001;
        16'b0000010011011010 : reciprocal = 16'b0000000000000001;
        16'b0000010011011011 : reciprocal = 16'b0000000000000001;
        16'b0000010011011100 : reciprocal = 16'b0000000000000001;
        16'b0000010011011101 : reciprocal = 16'b0000000000000001;
        16'b0000010011011110 : reciprocal = 16'b0000000000000001;
        16'b0000010011011111 : reciprocal = 16'b0000000000000001;
        16'b0000010011100000 : reciprocal = 16'b0000000000000001;
        16'b0000010011100001 : reciprocal = 16'b0000000000000001;
        16'b0000010011100010 : reciprocal = 16'b0000000000000001;
        16'b0000010011100011 : reciprocal = 16'b0000000000000001;
        16'b0000010011100100 : reciprocal = 16'b0000000000000001;
        16'b0000010011100101 : reciprocal = 16'b0000000000000001;
        16'b0000010011100110 : reciprocal = 16'b0000000000000001;
        16'b0000010011100111 : reciprocal = 16'b0000000000000001;
        16'b0000010011101000 : reciprocal = 16'b0000000000000001;
        16'b0000010011101001 : reciprocal = 16'b0000000000000001;
        16'b0000010011101010 : reciprocal = 16'b0000000000000001;
        16'b0000010011101011 : reciprocal = 16'b0000000000000001;
        16'b0000010011101100 : reciprocal = 16'b0000000000000001;
        16'b0000010011101101 : reciprocal = 16'b0000000000000001;
        16'b0000010011101110 : reciprocal = 16'b0000000000000001;
        16'b0000010011101111 : reciprocal = 16'b0000000000000001;
        16'b0000010011110000 : reciprocal = 16'b0000000000000001;
        16'b0000010011110001 : reciprocal = 16'b0000000000000001;
        16'b0000010011110010 : reciprocal = 16'b0000000000000001;
        16'b0000010011110011 : reciprocal = 16'b0000000000000001;
        16'b0000010011110100 : reciprocal = 16'b0000000000000001;
        16'b0000010011110101 : reciprocal = 16'b0000000000000001;
        16'b0000010011110110 : reciprocal = 16'b0000000000000001;
        16'b0000010011110111 : reciprocal = 16'b0000000000000001;
        16'b0000010011111000 : reciprocal = 16'b0000000000000001;
        16'b0000010011111001 : reciprocal = 16'b0000000000000001;
        16'b0000010011111010 : reciprocal = 16'b0000000000000001;
        16'b0000010011111011 : reciprocal = 16'b0000000000000001;
        16'b0000010011111100 : reciprocal = 16'b0000000000000001;
        16'b0000010011111101 : reciprocal = 16'b0000000000000001;
        16'b0000010011111110 : reciprocal = 16'b0000000000000001;
        16'b0000010011111111 : reciprocal = 16'b0000000000000001;
        16'b0000010100000000 : reciprocal = 16'b0000000000000001;
        16'b0000010100000001 : reciprocal = 16'b0000000000000001;
        16'b0000010100000010 : reciprocal = 16'b0000000000000001;
        16'b0000010100000011 : reciprocal = 16'b0000000000000001;
        16'b0000010100000100 : reciprocal = 16'b0000000000000001;
        16'b0000010100000101 : reciprocal = 16'b0000000000000001;
        16'b0000010100000110 : reciprocal = 16'b0000000000000001;
        16'b0000010100000111 : reciprocal = 16'b0000000000000001;
        16'b0000010100001000 : reciprocal = 16'b0000000000000001;
        16'b0000010100001001 : reciprocal = 16'b0000000000000001;
        16'b0000010100001010 : reciprocal = 16'b0000000000000001;
        16'b0000010100001011 : reciprocal = 16'b0000000000000001;
        16'b0000010100001100 : reciprocal = 16'b0000000000000001;
        16'b0000010100001101 : reciprocal = 16'b0000000000000001;
        16'b0000010100001110 : reciprocal = 16'b0000000000000001;
        16'b0000010100001111 : reciprocal = 16'b0000000000000001;
        16'b0000010100010000 : reciprocal = 16'b0000000000000001;
        16'b0000010100010001 : reciprocal = 16'b0000000000000001;
        16'b0000010100010010 : reciprocal = 16'b0000000000000001;
        16'b0000010100010011 : reciprocal = 16'b0000000000000001;
        16'b0000010100010100 : reciprocal = 16'b0000000000000001;
        16'b0000010100010101 : reciprocal = 16'b0000000000000001;
        16'b0000010100010110 : reciprocal = 16'b0000000000000001;
        16'b0000010100010111 : reciprocal = 16'b0000000000000001;
        16'b0000010100011000 : reciprocal = 16'b0000000000000001;
        16'b0000010100011001 : reciprocal = 16'b0000000000000001;
        16'b0000010100011010 : reciprocal = 16'b0000000000000001;
        16'b0000010100011011 : reciprocal = 16'b0000000000000001;
        16'b0000010100011100 : reciprocal = 16'b0000000000000001;
        16'b0000010100011101 : reciprocal = 16'b0000000000000001;
        16'b0000010100011110 : reciprocal = 16'b0000000000000001;
        16'b0000010100011111 : reciprocal = 16'b0000000000000001;
        16'b0000010100100000 : reciprocal = 16'b0000000000000001;
        16'b0000010100100001 : reciprocal = 16'b0000000000000001;
        16'b0000010100100010 : reciprocal = 16'b0000000000000001;
        16'b0000010100100011 : reciprocal = 16'b0000000000000001;
        16'b0000010100100100 : reciprocal = 16'b0000000000000001;
        16'b0000010100100101 : reciprocal = 16'b0000000000000001;
        16'b0000010100100110 : reciprocal = 16'b0000000000000001;
        16'b0000010100100111 : reciprocal = 16'b0000000000000001;
        16'b0000010100101000 : reciprocal = 16'b0000000000000001;
        16'b0000010100101001 : reciprocal = 16'b0000000000000001;
        16'b0000010100101010 : reciprocal = 16'b0000000000000001;
        16'b0000010100101011 : reciprocal = 16'b0000000000000001;
        16'b0000010100101100 : reciprocal = 16'b0000000000000001;
        16'b0000010100101101 : reciprocal = 16'b0000000000000001;
        16'b0000010100101110 : reciprocal = 16'b0000000000000001;
        16'b0000010100101111 : reciprocal = 16'b0000000000000001;
        16'b0000010100110000 : reciprocal = 16'b0000000000000001;
        16'b0000010100110001 : reciprocal = 16'b0000000000000001;
        16'b0000010100110010 : reciprocal = 16'b0000000000000001;
        16'b0000010100110011 : reciprocal = 16'b0000000000000001;
        16'b0000010100110100 : reciprocal = 16'b0000000000000001;
        16'b0000010100110101 : reciprocal = 16'b0000000000000001;
        16'b0000010100110110 : reciprocal = 16'b0000000000000001;
        16'b0000010100110111 : reciprocal = 16'b0000000000000001;
        16'b0000010100111000 : reciprocal = 16'b0000000000000001;
        16'b0000010100111001 : reciprocal = 16'b0000000000000001;
        16'b0000010100111010 : reciprocal = 16'b0000000000000001;
        16'b0000010100111011 : reciprocal = 16'b0000000000000001;
        16'b0000010100111100 : reciprocal = 16'b0000000000000001;
        16'b0000010100111101 : reciprocal = 16'b0000000000000001;
        16'b0000010100111110 : reciprocal = 16'b0000000000000001;
        16'b0000010100111111 : reciprocal = 16'b0000000000000001;
        16'b0000010101000000 : reciprocal = 16'b0000000000000001;
        16'b0000010101000001 : reciprocal = 16'b0000000000000001;
        16'b0000010101000010 : reciprocal = 16'b0000000000000001;
        16'b0000010101000011 : reciprocal = 16'b0000000000000001;
        16'b0000010101000100 : reciprocal = 16'b0000000000000001;
        16'b0000010101000101 : reciprocal = 16'b0000000000000001;
        16'b0000010101000110 : reciprocal = 16'b0000000000000001;
        16'b0000010101000111 : reciprocal = 16'b0000000000000001;
        16'b0000010101001000 : reciprocal = 16'b0000000000000001;
        16'b0000010101001001 : reciprocal = 16'b0000000000000001;
        16'b0000010101001010 : reciprocal = 16'b0000000000000001;
        16'b0000010101001011 : reciprocal = 16'b0000000000000001;
        16'b0000010101001100 : reciprocal = 16'b0000000000000001;
        16'b0000010101001101 : reciprocal = 16'b0000000000000001;
        16'b0000010101001110 : reciprocal = 16'b0000000000000001;
        16'b0000010101001111 : reciprocal = 16'b0000000000000001;
        16'b0000010101010000 : reciprocal = 16'b0000000000000001;
        16'b0000010101010001 : reciprocal = 16'b0000000000000001;
        16'b0000010101010010 : reciprocal = 16'b0000000000000001;
        16'b0000010101010011 : reciprocal = 16'b0000000000000001;
        16'b0000010101010100 : reciprocal = 16'b0000000000000001;
        16'b0000010101010101 : reciprocal = 16'b0000000000000001;
        16'b0000010101010110 : reciprocal = 16'b0000000000000001;
        16'b0000010101010111 : reciprocal = 16'b0000000000000001;
        16'b0000010101011000 : reciprocal = 16'b0000000000000001;
        16'b0000010101011001 : reciprocal = 16'b0000000000000001;
        16'b0000010101011010 : reciprocal = 16'b0000000000000001;
        16'b0000010101011011 : reciprocal = 16'b0000000000000001;
        16'b0000010101011100 : reciprocal = 16'b0000000000000001;
        16'b0000010101011101 : reciprocal = 16'b0000000000000001;
        16'b0000010101011110 : reciprocal = 16'b0000000000000001;
        16'b0000010101011111 : reciprocal = 16'b0000000000000001;
        16'b0000010101100000 : reciprocal = 16'b0000000000000001;
        16'b0000010101100001 : reciprocal = 16'b0000000000000001;
        16'b0000010101100010 : reciprocal = 16'b0000000000000001;
        16'b0000010101100011 : reciprocal = 16'b0000000000000001;
        16'b0000010101100100 : reciprocal = 16'b0000000000000001;
        16'b0000010101100101 : reciprocal = 16'b0000000000000001;
        16'b0000010101100110 : reciprocal = 16'b0000000000000001;
        16'b0000010101100111 : reciprocal = 16'b0000000000000001;
        16'b0000010101101000 : reciprocal = 16'b0000000000000001;
        16'b0000010101101001 : reciprocal = 16'b0000000000000001;
        16'b0000010101101010 : reciprocal = 16'b0000000000000001;
        16'b0000010101101011 : reciprocal = 16'b0000000000000001;
        16'b0000010101101100 : reciprocal = 16'b0000000000000001;
        16'b0000010101101101 : reciprocal = 16'b0000000000000001;
        16'b0000010101101110 : reciprocal = 16'b0000000000000001;
        16'b0000010101101111 : reciprocal = 16'b0000000000000001;
        16'b0000010101110000 : reciprocal = 16'b0000000000000001;
        16'b0000010101110001 : reciprocal = 16'b0000000000000001;
        16'b0000010101110010 : reciprocal = 16'b0000000000000001;
        16'b0000010101110011 : reciprocal = 16'b0000000000000001;
        16'b0000010101110100 : reciprocal = 16'b0000000000000001;
        16'b0000010101110101 : reciprocal = 16'b0000000000000001;
        16'b0000010101110110 : reciprocal = 16'b0000000000000001;
        16'b0000010101110111 : reciprocal = 16'b0000000000000001;
        16'b0000010101111000 : reciprocal = 16'b0000000000000001;
        16'b0000010101111001 : reciprocal = 16'b0000000000000001;
        16'b0000010101111010 : reciprocal = 16'b0000000000000001;
        16'b0000010101111011 : reciprocal = 16'b0000000000000001;
        16'b0000010101111100 : reciprocal = 16'b0000000000000001;
        16'b0000010101111101 : reciprocal = 16'b0000000000000001;
        16'b0000010101111110 : reciprocal = 16'b0000000000000001;
        16'b0000010101111111 : reciprocal = 16'b0000000000000001;
        16'b0000010110000000 : reciprocal = 16'b0000000000000001;
        16'b0000010110000001 : reciprocal = 16'b0000000000000001;
        16'b0000010110000010 : reciprocal = 16'b0000000000000001;
        16'b0000010110000011 : reciprocal = 16'b0000000000000001;
        16'b0000010110000100 : reciprocal = 16'b0000000000000001;
        16'b0000010110000101 : reciprocal = 16'b0000000000000001;
        16'b0000010110000110 : reciprocal = 16'b0000000000000001;
        16'b0000010110000111 : reciprocal = 16'b0000000000000001;
        16'b0000010110001000 : reciprocal = 16'b0000000000000001;
        16'b0000010110001001 : reciprocal = 16'b0000000000000001;
        16'b0000010110001010 : reciprocal = 16'b0000000000000001;
        16'b0000010110001011 : reciprocal = 16'b0000000000000001;
        16'b0000010110001100 : reciprocal = 16'b0000000000000001;
        16'b0000010110001101 : reciprocal = 16'b0000000000000001;
        16'b0000010110001110 : reciprocal = 16'b0000000000000001;
        16'b0000010110001111 : reciprocal = 16'b0000000000000001;
        16'b0000010110010000 : reciprocal = 16'b0000000000000001;
        16'b0000010110010001 : reciprocal = 16'b0000000000000001;
        16'b0000010110010010 : reciprocal = 16'b0000000000000001;
        16'b0000010110010011 : reciprocal = 16'b0000000000000001;
        16'b0000010110010100 : reciprocal = 16'b0000000000000001;
        16'b0000010110010101 : reciprocal = 16'b0000000000000001;
        16'b0000010110010110 : reciprocal = 16'b0000000000000001;
        16'b0000010110010111 : reciprocal = 16'b0000000000000001;
        16'b0000010110011000 : reciprocal = 16'b0000000000000001;
        16'b0000010110011001 : reciprocal = 16'b0000000000000001;
        16'b0000010110011010 : reciprocal = 16'b0000000000000001;
        16'b0000010110011011 : reciprocal = 16'b0000000000000001;
        16'b0000010110011100 : reciprocal = 16'b0000000000000001;
        16'b0000010110011101 : reciprocal = 16'b0000000000000001;
        16'b0000010110011110 : reciprocal = 16'b0000000000000001;
        16'b0000010110011111 : reciprocal = 16'b0000000000000001;
        16'b0000010110100000 : reciprocal = 16'b0000000000000001;
        16'b0000010110100001 : reciprocal = 16'b0000000000000001;
        16'b0000010110100010 : reciprocal = 16'b0000000000000001;
        16'b0000010110100011 : reciprocal = 16'b0000000000000001;
        16'b0000010110100100 : reciprocal = 16'b0000000000000001;
        16'b0000010110100101 : reciprocal = 16'b0000000000000001;
        16'b0000010110100110 : reciprocal = 16'b0000000000000001;
        16'b0000010110100111 : reciprocal = 16'b0000000000000001;
        16'b0000010110101000 : reciprocal = 16'b0000000000000001;
        16'b0000010110101001 : reciprocal = 16'b0000000000000001;
        16'b0000010110101010 : reciprocal = 16'b0000000000000001;
        16'b0000010110101011 : reciprocal = 16'b0000000000000001;
        16'b0000010110101100 : reciprocal = 16'b0000000000000001;
        16'b0000010110101101 : reciprocal = 16'b0000000000000001;
        16'b0000010110101110 : reciprocal = 16'b0000000000000001;
        16'b0000010110101111 : reciprocal = 16'b0000000000000001;
        16'b0000010110110000 : reciprocal = 16'b0000000000000001;
        16'b0000010110110001 : reciprocal = 16'b0000000000000001;
        16'b0000010110110010 : reciprocal = 16'b0000000000000001;
        16'b0000010110110011 : reciprocal = 16'b0000000000000001;
        16'b0000010110110100 : reciprocal = 16'b0000000000000001;
        16'b0000010110110101 : reciprocal = 16'b0000000000000001;
        16'b0000010110110110 : reciprocal = 16'b0000000000000001;
        16'b0000010110110111 : reciprocal = 16'b0000000000000001;
        16'b0000010110111000 : reciprocal = 16'b0000000000000001;
        16'b0000010110111001 : reciprocal = 16'b0000000000000001;
        16'b0000010110111010 : reciprocal = 16'b0000000000000001;
        16'b0000010110111011 : reciprocal = 16'b0000000000000001;
        16'b0000010110111100 : reciprocal = 16'b0000000000000001;
        16'b0000010110111101 : reciprocal = 16'b0000000000000001;
        16'b0000010110111110 : reciprocal = 16'b0000000000000001;
        16'b0000010110111111 : reciprocal = 16'b0000000000000001;
        16'b0000010111000000 : reciprocal = 16'b0000000000000001;
        16'b0000010111000001 : reciprocal = 16'b0000000000000001;
        16'b0000010111000010 : reciprocal = 16'b0000000000000001;
        16'b0000010111000011 : reciprocal = 16'b0000000000000001;
        16'b0000010111000100 : reciprocal = 16'b0000000000000001;
        16'b0000010111000101 : reciprocal = 16'b0000000000000001;
        16'b0000010111000110 : reciprocal = 16'b0000000000000001;
        16'b0000010111000111 : reciprocal = 16'b0000000000000001;
        16'b0000010111001000 : reciprocal = 16'b0000000000000001;
        16'b0000010111001001 : reciprocal = 16'b0000000000000001;
        16'b0000010111001010 : reciprocal = 16'b0000000000000001;
        16'b0000010111001011 : reciprocal = 16'b0000000000000001;
        16'b0000010111001100 : reciprocal = 16'b0000000000000001;
        16'b0000010111001101 : reciprocal = 16'b0000000000000001;
        16'b0000010111001110 : reciprocal = 16'b0000000000000001;
        16'b0000010111001111 : reciprocal = 16'b0000000000000001;
        16'b0000010111010000 : reciprocal = 16'b0000000000000001;
        16'b0000010111010001 : reciprocal = 16'b0000000000000001;
        16'b0000010111010010 : reciprocal = 16'b0000000000000001;
        16'b0000010111010011 : reciprocal = 16'b0000000000000001;
        16'b0000010111010100 : reciprocal = 16'b0000000000000001;
        16'b0000010111010101 : reciprocal = 16'b0000000000000001;
        16'b0000010111010110 : reciprocal = 16'b0000000000000001;
        16'b0000010111010111 : reciprocal = 16'b0000000000000001;
        16'b0000010111011000 : reciprocal = 16'b0000000000000001;
        16'b0000010111011001 : reciprocal = 16'b0000000000000001;
        16'b0000010111011010 : reciprocal = 16'b0000000000000001;
        16'b0000010111011011 : reciprocal = 16'b0000000000000001;
        16'b0000010111011100 : reciprocal = 16'b0000000000000001;
        16'b0000010111011101 : reciprocal = 16'b0000000000000001;
        16'b0000010111011110 : reciprocal = 16'b0000000000000001;
        16'b0000010111011111 : reciprocal = 16'b0000000000000001;
        16'b0000010111100000 : reciprocal = 16'b0000000000000001;
        16'b0000010111100001 : reciprocal = 16'b0000000000000001;
        16'b0000010111100010 : reciprocal = 16'b0000000000000001;
        16'b0000010111100011 : reciprocal = 16'b0000000000000001;
        16'b0000010111100100 : reciprocal = 16'b0000000000000001;
        16'b0000010111100101 : reciprocal = 16'b0000000000000001;
        16'b0000010111100110 : reciprocal = 16'b0000000000000001;
        16'b0000010111100111 : reciprocal = 16'b0000000000000001;
        16'b0000010111101000 : reciprocal = 16'b0000000000000001;
        16'b0000010111101001 : reciprocal = 16'b0000000000000001;
        16'b0000010111101010 : reciprocal = 16'b0000000000000001;
        16'b0000010111101011 : reciprocal = 16'b0000000000000001;
        16'b0000010111101100 : reciprocal = 16'b0000000000000001;
        16'b0000010111101101 : reciprocal = 16'b0000000000000001;
        16'b0000010111101110 : reciprocal = 16'b0000000000000001;
        16'b0000010111101111 : reciprocal = 16'b0000000000000001;
        16'b0000010111110000 : reciprocal = 16'b0000000000000001;
        16'b0000010111110001 : reciprocal = 16'b0000000000000001;
        16'b0000010111110010 : reciprocal = 16'b0000000000000001;
        16'b0000010111110011 : reciprocal = 16'b0000000000000001;
        16'b0000010111110100 : reciprocal = 16'b0000000000000001;
        16'b0000010111110101 : reciprocal = 16'b0000000000000001;
        16'b0000010111110110 : reciprocal = 16'b0000000000000001;
        16'b0000010111110111 : reciprocal = 16'b0000000000000001;
        16'b0000010111111000 : reciprocal = 16'b0000000000000001;
        16'b0000010111111001 : reciprocal = 16'b0000000000000001;
        16'b0000010111111010 : reciprocal = 16'b0000000000000001;
        16'b0000010111111011 : reciprocal = 16'b0000000000000001;
        16'b0000010111111100 : reciprocal = 16'b0000000000000001;
        16'b0000010111111101 : reciprocal = 16'b0000000000000001;
        16'b0000010111111110 : reciprocal = 16'b0000000000000001;
        16'b0000010111111111 : reciprocal = 16'b0000000000000001;
        16'b0000011000000000 : reciprocal = 16'b0000000000000001;
        16'b0000011000000001 : reciprocal = 16'b0000000000000001;
        16'b0000011000000010 : reciprocal = 16'b0000000000000001;
        16'b0000011000000011 : reciprocal = 16'b0000000000000001;
        16'b0000011000000100 : reciprocal = 16'b0000000000000001;
        16'b0000011000000101 : reciprocal = 16'b0000000000000001;
        16'b0000011000000110 : reciprocal = 16'b0000000000000001;
        16'b0000011000000111 : reciprocal = 16'b0000000000000001;
        16'b0000011000001000 : reciprocal = 16'b0000000000000001;
        16'b0000011000001001 : reciprocal = 16'b0000000000000001;
        16'b0000011000001010 : reciprocal = 16'b0000000000000001;
        16'b0000011000001011 : reciprocal = 16'b0000000000000001;
        16'b0000011000001100 : reciprocal = 16'b0000000000000001;
        16'b0000011000001101 : reciprocal = 16'b0000000000000001;
        16'b0000011000001110 : reciprocal = 16'b0000000000000001;
        16'b0000011000001111 : reciprocal = 16'b0000000000000001;
        16'b0000011000010000 : reciprocal = 16'b0000000000000001;
        16'b0000011000010001 : reciprocal = 16'b0000000000000001;
        16'b0000011000010010 : reciprocal = 16'b0000000000000001;
        16'b0000011000010011 : reciprocal = 16'b0000000000000001;
        16'b0000011000010100 : reciprocal = 16'b0000000000000001;
        16'b0000011000010101 : reciprocal = 16'b0000000000000001;
        16'b0000011000010110 : reciprocal = 16'b0000000000000001;
        16'b0000011000010111 : reciprocal = 16'b0000000000000001;
        16'b0000011000011000 : reciprocal = 16'b0000000000000001;
        16'b0000011000011001 : reciprocal = 16'b0000000000000001;
        16'b0000011000011010 : reciprocal = 16'b0000000000000001;
        16'b0000011000011011 : reciprocal = 16'b0000000000000001;
        16'b0000011000011100 : reciprocal = 16'b0000000000000001;
        16'b0000011000011101 : reciprocal = 16'b0000000000000001;
        16'b0000011000011110 : reciprocal = 16'b0000000000000001;
        16'b0000011000011111 : reciprocal = 16'b0000000000000001;
        16'b0000011000100000 : reciprocal = 16'b0000000000000001;
        16'b0000011000100001 : reciprocal = 16'b0000000000000001;
        16'b0000011000100010 : reciprocal = 16'b0000000000000001;
        16'b0000011000100011 : reciprocal = 16'b0000000000000001;
        16'b0000011000100100 : reciprocal = 16'b0000000000000001;
        16'b0000011000100101 : reciprocal = 16'b0000000000000001;
        16'b0000011000100110 : reciprocal = 16'b0000000000000001;
        16'b0000011000100111 : reciprocal = 16'b0000000000000001;
        16'b0000011000101000 : reciprocal = 16'b0000000000000001;
        16'b0000011000101001 : reciprocal = 16'b0000000000000001;
        16'b0000011000101010 : reciprocal = 16'b0000000000000001;
        16'b0000011000101011 : reciprocal = 16'b0000000000000001;
        16'b0000011000101100 : reciprocal = 16'b0000000000000001;
        16'b0000011000101101 : reciprocal = 16'b0000000000000001;
        16'b0000011000101110 : reciprocal = 16'b0000000000000001;
        16'b0000011000101111 : reciprocal = 16'b0000000000000001;
        16'b0000011000110000 : reciprocal = 16'b0000000000000001;
        16'b0000011000110001 : reciprocal = 16'b0000000000000001;
        16'b0000011000110010 : reciprocal = 16'b0000000000000001;
        16'b0000011000110011 : reciprocal = 16'b0000000000000001;
        16'b0000011000110100 : reciprocal = 16'b0000000000000001;
        16'b0000011000110101 : reciprocal = 16'b0000000000000001;
        16'b0000011000110110 : reciprocal = 16'b0000000000000001;
        16'b0000011000110111 : reciprocal = 16'b0000000000000001;
        16'b0000011000111000 : reciprocal = 16'b0000000000000001;
        16'b0000011000111001 : reciprocal = 16'b0000000000000001;
        16'b0000011000111010 : reciprocal = 16'b0000000000000001;
        16'b0000011000111011 : reciprocal = 16'b0000000000000001;
        16'b0000011000111100 : reciprocal = 16'b0000000000000001;
        16'b0000011000111101 : reciprocal = 16'b0000000000000001;
        16'b0000011000111110 : reciprocal = 16'b0000000000000001;
        16'b0000011000111111 : reciprocal = 16'b0000000000000001;
        16'b0000011001000000 : reciprocal = 16'b0000000000000001;
        16'b0000011001000001 : reciprocal = 16'b0000000000000001;
        16'b0000011001000010 : reciprocal = 16'b0000000000000001;
        16'b0000011001000011 : reciprocal = 16'b0000000000000001;
        16'b0000011001000100 : reciprocal = 16'b0000000000000001;
        16'b0000011001000101 : reciprocal = 16'b0000000000000001;
        16'b0000011001000110 : reciprocal = 16'b0000000000000001;
        16'b0000011001000111 : reciprocal = 16'b0000000000000001;
        16'b0000011001001000 : reciprocal = 16'b0000000000000001;
        16'b0000011001001001 : reciprocal = 16'b0000000000000001;
        16'b0000011001001010 : reciprocal = 16'b0000000000000001;
        16'b0000011001001011 : reciprocal = 16'b0000000000000001;
        16'b0000011001001100 : reciprocal = 16'b0000000000000001;
        16'b0000011001001101 : reciprocal = 16'b0000000000000001;
        16'b0000011001001110 : reciprocal = 16'b0000000000000001;
        16'b0000011001001111 : reciprocal = 16'b0000000000000001;
        16'b0000011001010000 : reciprocal = 16'b0000000000000001;
        16'b0000011001010001 : reciprocal = 16'b0000000000000001;
        16'b0000011001010010 : reciprocal = 16'b0000000000000001;
        16'b0000011001010011 : reciprocal = 16'b0000000000000001;
        16'b0000011001010100 : reciprocal = 16'b0000000000000001;
        16'b0000011001010101 : reciprocal = 16'b0000000000000001;
        16'b0000011001010110 : reciprocal = 16'b0000000000000001;
        16'b0000011001010111 : reciprocal = 16'b0000000000000001;
        16'b0000011001011000 : reciprocal = 16'b0000000000000001;
        16'b0000011001011001 : reciprocal = 16'b0000000000000001;
        16'b0000011001011010 : reciprocal = 16'b0000000000000001;
        16'b0000011001011011 : reciprocal = 16'b0000000000000001;
        16'b0000011001011100 : reciprocal = 16'b0000000000000001;
        16'b0000011001011101 : reciprocal = 16'b0000000000000001;
        16'b0000011001011110 : reciprocal = 16'b0000000000000001;
        16'b0000011001011111 : reciprocal = 16'b0000000000000001;
        16'b0000011001100000 : reciprocal = 16'b0000000000000001;
        16'b0000011001100001 : reciprocal = 16'b0000000000000001;
        16'b0000011001100010 : reciprocal = 16'b0000000000000001;
        16'b0000011001100011 : reciprocal = 16'b0000000000000001;
        16'b0000011001100100 : reciprocal = 16'b0000000000000001;
        16'b0000011001100101 : reciprocal = 16'b0000000000000001;
        16'b0000011001100110 : reciprocal = 16'b0000000000000001;
        16'b0000011001100111 : reciprocal = 16'b0000000000000001;
        16'b0000011001101000 : reciprocal = 16'b0000000000000001;
        16'b0000011001101001 : reciprocal = 16'b0000000000000001;
        16'b0000011001101010 : reciprocal = 16'b0000000000000001;
        16'b0000011001101011 : reciprocal = 16'b0000000000000001;
        16'b0000011001101100 : reciprocal = 16'b0000000000000001;
        16'b0000011001101101 : reciprocal = 16'b0000000000000001;
        16'b0000011001101110 : reciprocal = 16'b0000000000000001;
        16'b0000011001101111 : reciprocal = 16'b0000000000000001;
        16'b0000011001110000 : reciprocal = 16'b0000000000000001;
        16'b0000011001110001 : reciprocal = 16'b0000000000000001;
        16'b0000011001110010 : reciprocal = 16'b0000000000000001;
        16'b0000011001110011 : reciprocal = 16'b0000000000000001;
        16'b0000011001110100 : reciprocal = 16'b0000000000000001;
        16'b0000011001110101 : reciprocal = 16'b0000000000000001;
        16'b0000011001110110 : reciprocal = 16'b0000000000000001;
        16'b0000011001110111 : reciprocal = 16'b0000000000000001;
        16'b0000011001111000 : reciprocal = 16'b0000000000000001;
        16'b0000011001111001 : reciprocal = 16'b0000000000000001;
        16'b0000011001111010 : reciprocal = 16'b0000000000000001;
        16'b0000011001111011 : reciprocal = 16'b0000000000000001;
        16'b0000011001111100 : reciprocal = 16'b0000000000000001;
        16'b0000011001111101 : reciprocal = 16'b0000000000000001;
        16'b0000011001111110 : reciprocal = 16'b0000000000000001;
        16'b0000011001111111 : reciprocal = 16'b0000000000000001;
        16'b0000011010000000 : reciprocal = 16'b0000000000000001;
        16'b0000011010000001 : reciprocal = 16'b0000000000000001;
        16'b0000011010000010 : reciprocal = 16'b0000000000000001;
        16'b0000011010000011 : reciprocal = 16'b0000000000000001;
        16'b0000011010000100 : reciprocal = 16'b0000000000000001;
        16'b0000011010000101 : reciprocal = 16'b0000000000000001;
        16'b0000011010000110 : reciprocal = 16'b0000000000000001;
        16'b0000011010000111 : reciprocal = 16'b0000000000000001;
        16'b0000011010001000 : reciprocal = 16'b0000000000000001;
        16'b0000011010001001 : reciprocal = 16'b0000000000000001;
        16'b0000011010001010 : reciprocal = 16'b0000000000000001;
        16'b0000011010001011 : reciprocal = 16'b0000000000000001;
        16'b0000011010001100 : reciprocal = 16'b0000000000000001;
        16'b0000011010001101 : reciprocal = 16'b0000000000000001;
        16'b0000011010001110 : reciprocal = 16'b0000000000000001;
        16'b0000011010001111 : reciprocal = 16'b0000000000000001;
        16'b0000011010010000 : reciprocal = 16'b0000000000000001;
        16'b0000011010010001 : reciprocal = 16'b0000000000000001;
        16'b0000011010010010 : reciprocal = 16'b0000000000000001;
        16'b0000011010010011 : reciprocal = 16'b0000000000000001;
        16'b0000011010010100 : reciprocal = 16'b0000000000000001;
        16'b0000011010010101 : reciprocal = 16'b0000000000000001;
        16'b0000011010010110 : reciprocal = 16'b0000000000000001;
        16'b0000011010010111 : reciprocal = 16'b0000000000000001;
        16'b0000011010011000 : reciprocal = 16'b0000000000000001;
        16'b0000011010011001 : reciprocal = 16'b0000000000000001;
        16'b0000011010011010 : reciprocal = 16'b0000000000000001;
        16'b0000011010011011 : reciprocal = 16'b0000000000000001;
        16'b0000011010011100 : reciprocal = 16'b0000000000000001;
        16'b0000011010011101 : reciprocal = 16'b0000000000000001;
        16'b0000011010011110 : reciprocal = 16'b0000000000000001;
        16'b0000011010011111 : reciprocal = 16'b0000000000000001;
        16'b0000011010100000 : reciprocal = 16'b0000000000000001;
        16'b0000011010100001 : reciprocal = 16'b0000000000000001;
        16'b0000011010100010 : reciprocal = 16'b0000000000000001;
        16'b0000011010100011 : reciprocal = 16'b0000000000000001;
        16'b0000011010100100 : reciprocal = 16'b0000000000000001;
        16'b0000011010100101 : reciprocal = 16'b0000000000000001;
        16'b0000011010100110 : reciprocal = 16'b0000000000000001;
        16'b0000011010100111 : reciprocal = 16'b0000000000000001;
        16'b0000011010101000 : reciprocal = 16'b0000000000000001;
        16'b0000011010101001 : reciprocal = 16'b0000000000000001;
        16'b0000011010101010 : reciprocal = 16'b0000000000000001;
        16'b0000011010101011 : reciprocal = 16'b0000000000000001;
        16'b0000011010101100 : reciprocal = 16'b0000000000000001;
        16'b0000011010101101 : reciprocal = 16'b0000000000000001;
        16'b0000011010101110 : reciprocal = 16'b0000000000000001;
        16'b0000011010101111 : reciprocal = 16'b0000000000000001;
        16'b0000011010110000 : reciprocal = 16'b0000000000000001;
        16'b0000011010110001 : reciprocal = 16'b0000000000000001;
        16'b0000011010110010 : reciprocal = 16'b0000000000000001;
        16'b0000011010110011 : reciprocal = 16'b0000000000000001;
        16'b0000011010110100 : reciprocal = 16'b0000000000000001;
        16'b0000011010110101 : reciprocal = 16'b0000000000000001;
        16'b0000011010110110 : reciprocal = 16'b0000000000000001;
        16'b0000011010110111 : reciprocal = 16'b0000000000000001;
        16'b0000011010111000 : reciprocal = 16'b0000000000000001;
        16'b0000011010111001 : reciprocal = 16'b0000000000000001;
        16'b0000011010111010 : reciprocal = 16'b0000000000000001;
        16'b0000011010111011 : reciprocal = 16'b0000000000000001;
        16'b0000011010111100 : reciprocal = 16'b0000000000000001;
        16'b0000011010111101 : reciprocal = 16'b0000000000000001;
        16'b0000011010111110 : reciprocal = 16'b0000000000000001;
        16'b0000011010111111 : reciprocal = 16'b0000000000000001;
        16'b0000011011000000 : reciprocal = 16'b0000000000000001;
        16'b0000011011000001 : reciprocal = 16'b0000000000000001;
        16'b0000011011000010 : reciprocal = 16'b0000000000000001;
        16'b0000011011000011 : reciprocal = 16'b0000000000000001;
        16'b0000011011000100 : reciprocal = 16'b0000000000000001;
        16'b0000011011000101 : reciprocal = 16'b0000000000000001;
        16'b0000011011000110 : reciprocal = 16'b0000000000000001;
        16'b0000011011000111 : reciprocal = 16'b0000000000000001;
        16'b0000011011001000 : reciprocal = 16'b0000000000000001;
        16'b0000011011001001 : reciprocal = 16'b0000000000000001;
        16'b0000011011001010 : reciprocal = 16'b0000000000000001;
        16'b0000011011001011 : reciprocal = 16'b0000000000000001;
        16'b0000011011001100 : reciprocal = 16'b0000000000000001;
        16'b0000011011001101 : reciprocal = 16'b0000000000000001;
        16'b0000011011001110 : reciprocal = 16'b0000000000000001;
        16'b0000011011001111 : reciprocal = 16'b0000000000000001;
        16'b0000011011010000 : reciprocal = 16'b0000000000000001;
        16'b0000011011010001 : reciprocal = 16'b0000000000000001;
        16'b0000011011010010 : reciprocal = 16'b0000000000000001;
        16'b0000011011010011 : reciprocal = 16'b0000000000000001;
        16'b0000011011010100 : reciprocal = 16'b0000000000000001;
        16'b0000011011010101 : reciprocal = 16'b0000000000000001;
        16'b0000011011010110 : reciprocal = 16'b0000000000000001;
        16'b0000011011010111 : reciprocal = 16'b0000000000000001;
        16'b0000011011011000 : reciprocal = 16'b0000000000000001;
        16'b0000011011011001 : reciprocal = 16'b0000000000000001;
        16'b0000011011011010 : reciprocal = 16'b0000000000000001;
        16'b0000011011011011 : reciprocal = 16'b0000000000000001;
        16'b0000011011011100 : reciprocal = 16'b0000000000000001;
        16'b0000011011011101 : reciprocal = 16'b0000000000000001;
        16'b0000011011011110 : reciprocal = 16'b0000000000000001;
        16'b0000011011011111 : reciprocal = 16'b0000000000000001;
        16'b0000011011100000 : reciprocal = 16'b0000000000000001;
        16'b0000011011100001 : reciprocal = 16'b0000000000000001;
        16'b0000011011100010 : reciprocal = 16'b0000000000000001;
        16'b0000011011100011 : reciprocal = 16'b0000000000000001;
        16'b0000011011100100 : reciprocal = 16'b0000000000000001;
        16'b0000011011100101 : reciprocal = 16'b0000000000000001;
        16'b0000011011100110 : reciprocal = 16'b0000000000000001;
        16'b0000011011100111 : reciprocal = 16'b0000000000000001;
        16'b0000011011101000 : reciprocal = 16'b0000000000000001;
        16'b0000011011101001 : reciprocal = 16'b0000000000000001;
        16'b0000011011101010 : reciprocal = 16'b0000000000000001;
        16'b0000011011101011 : reciprocal = 16'b0000000000000001;
        16'b0000011011101100 : reciprocal = 16'b0000000000000001;
        16'b0000011011101101 : reciprocal = 16'b0000000000000001;
        16'b0000011011101110 : reciprocal = 16'b0000000000000001;
        16'b0000011011101111 : reciprocal = 16'b0000000000000001;
        16'b0000011011110000 : reciprocal = 16'b0000000000000001;
        16'b0000011011110001 : reciprocal = 16'b0000000000000001;
        16'b0000011011110010 : reciprocal = 16'b0000000000000001;
        16'b0000011011110011 : reciprocal = 16'b0000000000000001;
        16'b0000011011110100 : reciprocal = 16'b0000000000000001;
        16'b0000011011110101 : reciprocal = 16'b0000000000000001;
        16'b0000011011110110 : reciprocal = 16'b0000000000000001;
        16'b0000011011110111 : reciprocal = 16'b0000000000000001;
        16'b0000011011111000 : reciprocal = 16'b0000000000000001;
        16'b0000011011111001 : reciprocal = 16'b0000000000000001;
        16'b0000011011111010 : reciprocal = 16'b0000000000000001;
        16'b0000011011111011 : reciprocal = 16'b0000000000000001;
        16'b0000011011111100 : reciprocal = 16'b0000000000000001;
        16'b0000011011111101 : reciprocal = 16'b0000000000000001;
        16'b0000011011111110 : reciprocal = 16'b0000000000000001;
        16'b0000011011111111 : reciprocal = 16'b0000000000000001;
        16'b0000011100000000 : reciprocal = 16'b0000000000000001;
        16'b0000011100000001 : reciprocal = 16'b0000000000000001;
        16'b0000011100000010 : reciprocal = 16'b0000000000000001;
        16'b0000011100000011 : reciprocal = 16'b0000000000000001;
        16'b0000011100000100 : reciprocal = 16'b0000000000000001;
        16'b0000011100000101 : reciprocal = 16'b0000000000000001;
        16'b0000011100000110 : reciprocal = 16'b0000000000000001;
        16'b0000011100000111 : reciprocal = 16'b0000000000000001;
        16'b0000011100001000 : reciprocal = 16'b0000000000000001;
        16'b0000011100001001 : reciprocal = 16'b0000000000000001;
        16'b0000011100001010 : reciprocal = 16'b0000000000000001;
        16'b0000011100001011 : reciprocal = 16'b0000000000000001;
        16'b0000011100001100 : reciprocal = 16'b0000000000000001;
        16'b0000011100001101 : reciprocal = 16'b0000000000000001;
        16'b0000011100001110 : reciprocal = 16'b0000000000000001;
        16'b0000011100001111 : reciprocal = 16'b0000000000000001;
        16'b0000011100010000 : reciprocal = 16'b0000000000000001;
        16'b0000011100010001 : reciprocal = 16'b0000000000000001;
        16'b0000011100010010 : reciprocal = 16'b0000000000000001;
        16'b0000011100010011 : reciprocal = 16'b0000000000000001;
        16'b0000011100010100 : reciprocal = 16'b0000000000000001;
        16'b0000011100010101 : reciprocal = 16'b0000000000000001;
        16'b0000011100010110 : reciprocal = 16'b0000000000000001;
        16'b0000011100010111 : reciprocal = 16'b0000000000000001;
        16'b0000011100011000 : reciprocal = 16'b0000000000000001;
        16'b0000011100011001 : reciprocal = 16'b0000000000000001;
        16'b0000011100011010 : reciprocal = 16'b0000000000000001;
        16'b0000011100011011 : reciprocal = 16'b0000000000000001;
        16'b0000011100011100 : reciprocal = 16'b0000000000000001;
        16'b0000011100011101 : reciprocal = 16'b0000000000000001;
        16'b0000011100011110 : reciprocal = 16'b0000000000000001;
        16'b0000011100011111 : reciprocal = 16'b0000000000000001;
        16'b0000011100100000 : reciprocal = 16'b0000000000000001;
        16'b0000011100100001 : reciprocal = 16'b0000000000000001;
        16'b0000011100100010 : reciprocal = 16'b0000000000000001;
        16'b0000011100100011 : reciprocal = 16'b0000000000000001;
        16'b0000011100100100 : reciprocal = 16'b0000000000000001;
        16'b0000011100100101 : reciprocal = 16'b0000000000000001;
        16'b0000011100100110 : reciprocal = 16'b0000000000000001;
        16'b0000011100100111 : reciprocal = 16'b0000000000000001;
        16'b0000011100101000 : reciprocal = 16'b0000000000000001;
        16'b0000011100101001 : reciprocal = 16'b0000000000000001;
        16'b0000011100101010 : reciprocal = 16'b0000000000000001;
        16'b0000011100101011 : reciprocal = 16'b0000000000000001;
        16'b0000011100101100 : reciprocal = 16'b0000000000000001;
        16'b0000011100101101 : reciprocal = 16'b0000000000000001;
        16'b0000011100101110 : reciprocal = 16'b0000000000000001;
        16'b0000011100101111 : reciprocal = 16'b0000000000000001;
        16'b0000011100110000 : reciprocal = 16'b0000000000000001;
        16'b0000011100110001 : reciprocal = 16'b0000000000000001;
        16'b0000011100110010 : reciprocal = 16'b0000000000000001;
        16'b0000011100110011 : reciprocal = 16'b0000000000000001;
        16'b0000011100110100 : reciprocal = 16'b0000000000000001;
        16'b0000011100110101 : reciprocal = 16'b0000000000000001;
        16'b0000011100110110 : reciprocal = 16'b0000000000000001;
        16'b0000011100110111 : reciprocal = 16'b0000000000000001;
        16'b0000011100111000 : reciprocal = 16'b0000000000000001;
        16'b0000011100111001 : reciprocal = 16'b0000000000000001;
        16'b0000011100111010 : reciprocal = 16'b0000000000000001;
        16'b0000011100111011 : reciprocal = 16'b0000000000000001;
        16'b0000011100111100 : reciprocal = 16'b0000000000000001;
        16'b0000011100111101 : reciprocal = 16'b0000000000000001;
        16'b0000011100111110 : reciprocal = 16'b0000000000000001;
        16'b0000011100111111 : reciprocal = 16'b0000000000000001;
        16'b0000011101000000 : reciprocal = 16'b0000000000000001;
        16'b0000011101000001 : reciprocal = 16'b0000000000000001;
        16'b0000011101000010 : reciprocal = 16'b0000000000000001;
        16'b0000011101000011 : reciprocal = 16'b0000000000000001;
        16'b0000011101000100 : reciprocal = 16'b0000000000000001;
        16'b0000011101000101 : reciprocal = 16'b0000000000000001;
        16'b0000011101000110 : reciprocal = 16'b0000000000000001;
        16'b0000011101000111 : reciprocal = 16'b0000000000000001;
        16'b0000011101001000 : reciprocal = 16'b0000000000000001;
        16'b0000011101001001 : reciprocal = 16'b0000000000000001;
        16'b0000011101001010 : reciprocal = 16'b0000000000000001;
        16'b0000011101001011 : reciprocal = 16'b0000000000000001;
        16'b0000011101001100 : reciprocal = 16'b0000000000000001;
        16'b0000011101001101 : reciprocal = 16'b0000000000000001;
        16'b0000011101001110 : reciprocal = 16'b0000000000000001;
        16'b0000011101001111 : reciprocal = 16'b0000000000000001;
        16'b0000011101010000 : reciprocal = 16'b0000000000000001;
        16'b0000011101010001 : reciprocal = 16'b0000000000000001;
        16'b0000011101010010 : reciprocal = 16'b0000000000000001;
        16'b0000011101010011 : reciprocal = 16'b0000000000000001;
        16'b0000011101010100 : reciprocal = 16'b0000000000000001;
        16'b0000011101010101 : reciprocal = 16'b0000000000000001;
        16'b0000011101010110 : reciprocal = 16'b0000000000000001;
        16'b0000011101010111 : reciprocal = 16'b0000000000000001;
        16'b0000011101011000 : reciprocal = 16'b0000000000000001;
        16'b0000011101011001 : reciprocal = 16'b0000000000000001;
        16'b0000011101011010 : reciprocal = 16'b0000000000000001;
        16'b0000011101011011 : reciprocal = 16'b0000000000000001;
        16'b0000011101011100 : reciprocal = 16'b0000000000000001;
        16'b0000011101011101 : reciprocal = 16'b0000000000000001;
        16'b0000011101011110 : reciprocal = 16'b0000000000000001;
        16'b0000011101011111 : reciprocal = 16'b0000000000000001;
        16'b0000011101100000 : reciprocal = 16'b0000000000000001;
        16'b0000011101100001 : reciprocal = 16'b0000000000000001;
        16'b0000011101100010 : reciprocal = 16'b0000000000000001;
        16'b0000011101100011 : reciprocal = 16'b0000000000000001;
        16'b0000011101100100 : reciprocal = 16'b0000000000000001;
        16'b0000011101100101 : reciprocal = 16'b0000000000000001;
        16'b0000011101100110 : reciprocal = 16'b0000000000000001;
        16'b0000011101100111 : reciprocal = 16'b0000000000000001;
        16'b0000011101101000 : reciprocal = 16'b0000000000000001;
        16'b0000011101101001 : reciprocal = 16'b0000000000000001;
        16'b0000011101101010 : reciprocal = 16'b0000000000000001;
        16'b0000011101101011 : reciprocal = 16'b0000000000000001;
        16'b0000011101101100 : reciprocal = 16'b0000000000000001;
        16'b0000011101101101 : reciprocal = 16'b0000000000000001;
        16'b0000011101101110 : reciprocal = 16'b0000000000000001;
        16'b0000011101101111 : reciprocal = 16'b0000000000000001;
        16'b0000011101110000 : reciprocal = 16'b0000000000000001;
        16'b0000011101110001 : reciprocal = 16'b0000000000000001;
        16'b0000011101110010 : reciprocal = 16'b0000000000000001;
        16'b0000011101110011 : reciprocal = 16'b0000000000000001;
        16'b0000011101110100 : reciprocal = 16'b0000000000000001;
        16'b0000011101110101 : reciprocal = 16'b0000000000000001;
        16'b0000011101110110 : reciprocal = 16'b0000000000000001;
        16'b0000011101110111 : reciprocal = 16'b0000000000000001;
        16'b0000011101111000 : reciprocal = 16'b0000000000000001;
        16'b0000011101111001 : reciprocal = 16'b0000000000000001;
        16'b0000011101111010 : reciprocal = 16'b0000000000000001;
        16'b0000011101111011 : reciprocal = 16'b0000000000000001;
        16'b0000011101111100 : reciprocal = 16'b0000000000000001;
        16'b0000011101111101 : reciprocal = 16'b0000000000000001;
        16'b0000011101111110 : reciprocal = 16'b0000000000000001;
        16'b0000011101111111 : reciprocal = 16'b0000000000000001;
        16'b0000011110000000 : reciprocal = 16'b0000000000000001;
        16'b0000011110000001 : reciprocal = 16'b0000000000000001;
        16'b0000011110000010 : reciprocal = 16'b0000000000000001;
        16'b0000011110000011 : reciprocal = 16'b0000000000000001;
        16'b0000011110000100 : reciprocal = 16'b0000000000000001;
        16'b0000011110000101 : reciprocal = 16'b0000000000000001;
        16'b0000011110000110 : reciprocal = 16'b0000000000000001;
        16'b0000011110000111 : reciprocal = 16'b0000000000000001;
        16'b0000011110001000 : reciprocal = 16'b0000000000000001;
        16'b0000011110001001 : reciprocal = 16'b0000000000000001;
        16'b0000011110001010 : reciprocal = 16'b0000000000000001;
        16'b0000011110001011 : reciprocal = 16'b0000000000000001;
        16'b0000011110001100 : reciprocal = 16'b0000000000000001;
        16'b0000011110001101 : reciprocal = 16'b0000000000000001;
        16'b0000011110001110 : reciprocal = 16'b0000000000000001;
        16'b0000011110001111 : reciprocal = 16'b0000000000000001;
        16'b0000011110010000 : reciprocal = 16'b0000000000000001;
        16'b0000011110010001 : reciprocal = 16'b0000000000000001;
        16'b0000011110010010 : reciprocal = 16'b0000000000000001;
        16'b0000011110010011 : reciprocal = 16'b0000000000000001;
        16'b0000011110010100 : reciprocal = 16'b0000000000000001;
        16'b0000011110010101 : reciprocal = 16'b0000000000000001;
        16'b0000011110010110 : reciprocal = 16'b0000000000000001;
        16'b0000011110010111 : reciprocal = 16'b0000000000000001;
        16'b0000011110011000 : reciprocal = 16'b0000000000000001;
        16'b0000011110011001 : reciprocal = 16'b0000000000000001;
        16'b0000011110011010 : reciprocal = 16'b0000000000000001;
        16'b0000011110011011 : reciprocal = 16'b0000000000000001;
        16'b0000011110011100 : reciprocal = 16'b0000000000000001;
        16'b0000011110011101 : reciprocal = 16'b0000000000000001;
        16'b0000011110011110 : reciprocal = 16'b0000000000000001;
        16'b0000011110011111 : reciprocal = 16'b0000000000000001;
        16'b0000011110100000 : reciprocal = 16'b0000000000000001;
        16'b0000011110100001 : reciprocal = 16'b0000000000000001;
        16'b0000011110100010 : reciprocal = 16'b0000000000000001;
        16'b0000011110100011 : reciprocal = 16'b0000000000000001;
        16'b0000011110100100 : reciprocal = 16'b0000000000000001;
        16'b0000011110100101 : reciprocal = 16'b0000000000000001;
        16'b0000011110100110 : reciprocal = 16'b0000000000000001;
        16'b0000011110100111 : reciprocal = 16'b0000000000000001;
        16'b0000011110101000 : reciprocal = 16'b0000000000000001;
        16'b0000011110101001 : reciprocal = 16'b0000000000000001;
        16'b0000011110101010 : reciprocal = 16'b0000000000000001;
        16'b0000011110101011 : reciprocal = 16'b0000000000000001;
        16'b0000011110101100 : reciprocal = 16'b0000000000000001;
        16'b0000011110101101 : reciprocal = 16'b0000000000000001;
        16'b0000011110101110 : reciprocal = 16'b0000000000000001;
        16'b0000011110101111 : reciprocal = 16'b0000000000000001;
        16'b0000011110110000 : reciprocal = 16'b0000000000000001;
        16'b0000011110110001 : reciprocal = 16'b0000000000000001;
        16'b0000011110110010 : reciprocal = 16'b0000000000000001;
        16'b0000011110110011 : reciprocal = 16'b0000000000000001;
        16'b0000011110110100 : reciprocal = 16'b0000000000000001;
        16'b0000011110110101 : reciprocal = 16'b0000000000000001;
        16'b0000011110110110 : reciprocal = 16'b0000000000000001;
        16'b0000011110110111 : reciprocal = 16'b0000000000000001;
        16'b0000011110111000 : reciprocal = 16'b0000000000000001;
        16'b0000011110111001 : reciprocal = 16'b0000000000000001;
        16'b0000011110111010 : reciprocal = 16'b0000000000000001;
        16'b0000011110111011 : reciprocal = 16'b0000000000000001;
        16'b0000011110111100 : reciprocal = 16'b0000000000000001;
        16'b0000011110111101 : reciprocal = 16'b0000000000000001;
        16'b0000011110111110 : reciprocal = 16'b0000000000000001;
        16'b0000011110111111 : reciprocal = 16'b0000000000000001;
        16'b0000011111000000 : reciprocal = 16'b0000000000000001;
        16'b0000011111000001 : reciprocal = 16'b0000000000000001;
        16'b0000011111000010 : reciprocal = 16'b0000000000000001;
        16'b0000011111000011 : reciprocal = 16'b0000000000000001;
        16'b0000011111000100 : reciprocal = 16'b0000000000000001;
        16'b0000011111000101 : reciprocal = 16'b0000000000000001;
        16'b0000011111000110 : reciprocal = 16'b0000000000000001;
        16'b0000011111000111 : reciprocal = 16'b0000000000000001;
        16'b0000011111001000 : reciprocal = 16'b0000000000000001;
        16'b0000011111001001 : reciprocal = 16'b0000000000000001;
        16'b0000011111001010 : reciprocal = 16'b0000000000000001;
        16'b0000011111001011 : reciprocal = 16'b0000000000000001;
        16'b0000011111001100 : reciprocal = 16'b0000000000000001;
        16'b0000011111001101 : reciprocal = 16'b0000000000000001;
        16'b0000011111001110 : reciprocal = 16'b0000000000000001;
        16'b0000011111001111 : reciprocal = 16'b0000000000000001;
        16'b0000011111010000 : reciprocal = 16'b0000000000000001;
        16'b0000011111010001 : reciprocal = 16'b0000000000000001;
        16'b0000011111010010 : reciprocal = 16'b0000000000000001;
        16'b0000011111010011 : reciprocal = 16'b0000000000000001;
        16'b0000011111010100 : reciprocal = 16'b0000000000000001;
        16'b0000011111010101 : reciprocal = 16'b0000000000000001;
        16'b0000011111010110 : reciprocal = 16'b0000000000000001;
        16'b0000011111010111 : reciprocal = 16'b0000000000000001;
        16'b0000011111011000 : reciprocal = 16'b0000000000000001;
        16'b0000011111011001 : reciprocal = 16'b0000000000000001;
        16'b0000011111011010 : reciprocal = 16'b0000000000000001;
        16'b0000011111011011 : reciprocal = 16'b0000000000000001;
        16'b0000011111011100 : reciprocal = 16'b0000000000000001;
        16'b0000011111011101 : reciprocal = 16'b0000000000000001;
        16'b0000011111011110 : reciprocal = 16'b0000000000000001;
        16'b0000011111011111 : reciprocal = 16'b0000000000000001;
        16'b0000011111100000 : reciprocal = 16'b0000000000000001;
        16'b0000011111100001 : reciprocal = 16'b0000000000000001;
        16'b0000011111100010 : reciprocal = 16'b0000000000000001;
        16'b0000011111100011 : reciprocal = 16'b0000000000000001;
        16'b0000011111100100 : reciprocal = 16'b0000000000000001;
        16'b0000011111100101 : reciprocal = 16'b0000000000000001;
        16'b0000011111100110 : reciprocal = 16'b0000000000000001;
        16'b0000011111100111 : reciprocal = 16'b0000000000000001;
        16'b0000011111101000 : reciprocal = 16'b0000000000000001;
        16'b0000011111101001 : reciprocal = 16'b0000000000000001;
        16'b0000011111101010 : reciprocal = 16'b0000000000000001;
        16'b0000011111101011 : reciprocal = 16'b0000000000000001;
        16'b0000011111101100 : reciprocal = 16'b0000000000000001;
        16'b0000011111101101 : reciprocal = 16'b0000000000000001;
        16'b0000011111101110 : reciprocal = 16'b0000000000000001;
        16'b0000011111101111 : reciprocal = 16'b0000000000000001;
        16'b0000011111110000 : reciprocal = 16'b0000000000000001;
        16'b0000011111110001 : reciprocal = 16'b0000000000000001;
        16'b0000011111110010 : reciprocal = 16'b0000000000000001;
        16'b0000011111110011 : reciprocal = 16'b0000000000000001;
        16'b0000011111110100 : reciprocal = 16'b0000000000000001;
        16'b0000011111110101 : reciprocal = 16'b0000000000000001;
        16'b0000011111110110 : reciprocal = 16'b0000000000000001;
        16'b0000011111110111 : reciprocal = 16'b0000000000000001;
        16'b0000011111111000 : reciprocal = 16'b0000000000000001;
        16'b0000011111111001 : reciprocal = 16'b0000000000000001;
        16'b0000011111111010 : reciprocal = 16'b0000000000000001;
        16'b0000011111111011 : reciprocal = 16'b0000000000000001;
        16'b0000011111111100 : reciprocal = 16'b0000000000000001;
        16'b0000011111111101 : reciprocal = 16'b0000000000000001;
        16'b0000011111111110 : reciprocal = 16'b0000000000000001;
        16'b0000011111111111 : reciprocal = 16'b0000000000000001;
        default : reciprocal = 16'b0000000000000000;
        16'b1111111111111111 : reciprocal = 1111110000000000;
        16'b1111111111111110 : reciprocal = 1111111000000000;
        16'b1111111111111101 : reciprocal = 1111111010101011;
        16'b1111111111111100 : reciprocal = 1111111100000000;
        16'b1111111111111011 : reciprocal = 1111111100110011;
        16'b1111111111111010 : reciprocal = 1111111101010101;
        16'b1111111111111001 : reciprocal = 1111111101101110;
        16'b1111111111111000 : reciprocal = 1111111110000000;
        16'b1111111111110111 : reciprocal = 1111111110001110;
        16'b1111111111110110 : reciprocal = 1111111110011010;
        16'b1111111111110101 : reciprocal = 1111111110100011;
        16'b1111111111110100 : reciprocal = 1111111110101011;
        16'b1111111111110011 : reciprocal = 1111111110110001;
        16'b1111111111110010 : reciprocal = 1111111110110111;
        16'b1111111111110001 : reciprocal = 1111111110111100;
        16'b1111111111110000 : reciprocal = 1111111111000000;
        16'b1111111111101111 : reciprocal = 1111111111000100;
        16'b1111111111101110 : reciprocal = 1111111111000111;
        16'b1111111111101101 : reciprocal = 1111111111001010;
        16'b1111111111101100 : reciprocal = 1111111111001101;
        16'b1111111111101011 : reciprocal = 1111111111001111;
        16'b1111111111101010 : reciprocal = 1111111111010001;
        16'b1111111111101001 : reciprocal = 1111111111010011;
        16'b1111111111101000 : reciprocal = 1111111111010101;
        16'b1111111111100111 : reciprocal = 1111111111010111;
        16'b1111111111100110 : reciprocal = 1111111111011001;
        16'b1111111111100101 : reciprocal = 1111111111011010;
        16'b1111111111100100 : reciprocal = 1111111111011011;
        16'b1111111111100011 : reciprocal = 1111111111011101;
        16'b1111111111100010 : reciprocal = 1111111111011110;
        16'b1111111111100001 : reciprocal = 1111111111011111;
        16'b1111111111100000 : reciprocal = 1111111111100000;
        16'b1111111111011111 : reciprocal = 1111111111100001;
        16'b1111111111011110 : reciprocal = 1111111111100010;
        16'b1111111111011101 : reciprocal = 1111111111100011;
        16'b1111111111011100 : reciprocal = 1111111111100100;
        16'b1111111111011011 : reciprocal = 1111111111100100;
        16'b1111111111011010 : reciprocal = 1111111111100101;
        16'b1111111111011001 : reciprocal = 1111111111100110;
        16'b1111111111011000 : reciprocal = 1111111111100110;
        16'b1111111111010111 : reciprocal = 1111111111100111;
        16'b1111111111010110 : reciprocal = 1111111111101000;
        16'b1111111111010101 : reciprocal = 1111111111101000;
        16'b1111111111010100 : reciprocal = 1111111111101001;
        16'b1111111111010011 : reciprocal = 1111111111101001;
        16'b1111111111010010 : reciprocal = 1111111111101010;
        16'b1111111111010001 : reciprocal = 1111111111101010;
        16'b1111111111010000 : reciprocal = 1111111111101011;
        16'b1111111111001111 : reciprocal = 1111111111101011;
        16'b1111111111001110 : reciprocal = 1111111111101100;
        16'b1111111111001101 : reciprocal = 1111111111101100;
        16'b1111111111001100 : reciprocal = 1111111111101100;
        16'b1111111111001011 : reciprocal = 1111111111101101;
        16'b1111111111001010 : reciprocal = 1111111111101101;
        16'b1111111111001001 : reciprocal = 1111111111101101;
        16'b1111111111001000 : reciprocal = 1111111111101110;
        16'b1111111111000111 : reciprocal = 1111111111101110;
        16'b1111111111000110 : reciprocal = 1111111111101110;
        16'b1111111111000101 : reciprocal = 1111111111101111;
        16'b1111111111000100 : reciprocal = 1111111111101111;
        16'b1111111111000011 : reciprocal = 1111111111101111;
        16'b1111111111000010 : reciprocal = 1111111111101111;
        16'b1111111111000001 : reciprocal = 1111111111110000;
        16'b1111111111000000 : reciprocal = 1111111111110000;
        16'b1111111110111111 : reciprocal = 1111111111110000;
        16'b1111111110111110 : reciprocal = 1111111111110000;
        16'b1111111110111101 : reciprocal = 1111111111110001;
        16'b1111111110111100 : reciprocal = 1111111111110001;
        16'b1111111110111011 : reciprocal = 1111111111110001;
        16'b1111111110111010 : reciprocal = 1111111111110001;
        16'b1111111110111001 : reciprocal = 1111111111110010;
        16'b1111111110111000 : reciprocal = 1111111111110010;
        16'b1111111110110111 : reciprocal = 1111111111110010;
        16'b1111111110110110 : reciprocal = 1111111111110010;
        16'b1111111110110101 : reciprocal = 1111111111110010;
        16'b1111111110110100 : reciprocal = 1111111111110011;
        16'b1111111110110011 : reciprocal = 1111111111110011;
        16'b1111111110110010 : reciprocal = 1111111111110011;
        16'b1111111110110001 : reciprocal = 1111111111110011;
        16'b1111111110110000 : reciprocal = 1111111111110011;
        16'b1111111110101111 : reciprocal = 1111111111110011;
        16'b1111111110101110 : reciprocal = 1111111111110100;
        16'b1111111110101101 : reciprocal = 1111111111110100;
        16'b1111111110101100 : reciprocal = 1111111111110100;
        16'b1111111110101011 : reciprocal = 1111111111110100;
        16'b1111111110101010 : reciprocal = 1111111111110100;
        16'b1111111110101001 : reciprocal = 1111111111110100;
        16'b1111111110101000 : reciprocal = 1111111111110100;
        16'b1111111110100111 : reciprocal = 1111111111110100;
        16'b1111111110100110 : reciprocal = 1111111111110101;
        16'b1111111110100101 : reciprocal = 1111111111110101;
        16'b1111111110100100 : reciprocal = 1111111111110101;
        16'b1111111110100011 : reciprocal = 1111111111110101;
        16'b1111111110100010 : reciprocal = 1111111111110101;
        16'b1111111110100001 : reciprocal = 1111111111110101;
        16'b1111111110100000 : reciprocal = 1111111111110101;
        16'b1111111110011111 : reciprocal = 1111111111110101;
        16'b1111111110011110 : reciprocal = 1111111111110110;
        16'b1111111110011101 : reciprocal = 1111111111110110;
        16'b1111111110011100 : reciprocal = 1111111111110110;
        16'b1111111110011011 : reciprocal = 1111111111110110;
        16'b1111111110011010 : reciprocal = 1111111111110110;
        16'b1111111110011001 : reciprocal = 1111111111110110;
        16'b1111111110011000 : reciprocal = 1111111111110110;
        16'b1111111110010111 : reciprocal = 1111111111110110;
        16'b1111111110010110 : reciprocal = 1111111111110110;
        16'b1111111110010101 : reciprocal = 1111111111110110;
        16'b1111111110010100 : reciprocal = 1111111111110111;
        16'b1111111110010011 : reciprocal = 1111111111110111;
        16'b1111111110010010 : reciprocal = 1111111111110111;
        16'b1111111110010001 : reciprocal = 1111111111110111;
        16'b1111111110010000 : reciprocal = 1111111111110111;
        16'b1111111110001111 : reciprocal = 1111111111110111;
        16'b1111111110001110 : reciprocal = 1111111111110111;
        16'b1111111110001101 : reciprocal = 1111111111110111;
        16'b1111111110001100 : reciprocal = 1111111111110111;
        16'b1111111110001011 : reciprocal = 1111111111110111;
        16'b1111111110001010 : reciprocal = 1111111111110111;
        16'b1111111110001001 : reciprocal = 1111111111110111;
        16'b1111111110001000 : reciprocal = 1111111111110111;
        16'b1111111110000111 : reciprocal = 1111111111111000;
        16'b1111111110000110 : reciprocal = 1111111111111000;
        16'b1111111110000101 : reciprocal = 1111111111111000;
        16'b1111111110000100 : reciprocal = 1111111111111000;
        16'b1111111110000011 : reciprocal = 1111111111111000;
        16'b1111111110000010 : reciprocal = 1111111111111000;
        16'b1111111110000001 : reciprocal = 1111111111111000;
        16'b1111111110000000 : reciprocal = 1111111111111000;
        16'b1111111101111111 : reciprocal = 1111111111111000;
        16'b1111111101111110 : reciprocal = 1111111111111000;
        16'b1111111101111101 : reciprocal = 1111111111111000;
        16'b1111111101111100 : reciprocal = 1111111111111000;
        16'b1111111101111011 : reciprocal = 1111111111111000;
        16'b1111111101111010 : reciprocal = 1111111111111000;
        16'b1111111101111001 : reciprocal = 1111111111111000;
        16'b1111111101111000 : reciprocal = 1111111111111000;
        16'b1111111101110111 : reciprocal = 1111111111111001;
        16'b1111111101110110 : reciprocal = 1111111111111001;
        16'b1111111101110101 : reciprocal = 1111111111111001;
        16'b1111111101110100 : reciprocal = 1111111111111001;
        16'b1111111101110011 : reciprocal = 1111111111111001;
        16'b1111111101110010 : reciprocal = 1111111111111001;
        16'b1111111101110001 : reciprocal = 1111111111111001;
        16'b1111111101110000 : reciprocal = 1111111111111001;
        16'b1111111101101111 : reciprocal = 1111111111111001;
        16'b1111111101101110 : reciprocal = 1111111111111001;
        16'b1111111101101101 : reciprocal = 1111111111111001;
        16'b1111111101101100 : reciprocal = 1111111111111001;
        16'b1111111101101011 : reciprocal = 1111111111111001;
        16'b1111111101101010 : reciprocal = 1111111111111001;
        16'b1111111101101001 : reciprocal = 1111111111111001;
        16'b1111111101101000 : reciprocal = 1111111111111001;
        16'b1111111101100111 : reciprocal = 1111111111111001;
        16'b1111111101100110 : reciprocal = 1111111111111001;
        16'b1111111101100101 : reciprocal = 1111111111111001;
        16'b1111111101100100 : reciprocal = 1111111111111001;
        16'b1111111101100011 : reciprocal = 1111111111111001;
        16'b1111111101100010 : reciprocal = 1111111111111010;
        16'b1111111101100001 : reciprocal = 1111111111111010;
        16'b1111111101100000 : reciprocal = 1111111111111010;
        16'b1111111101011111 : reciprocal = 1111111111111010;
        16'b1111111101011110 : reciprocal = 1111111111111010;
        16'b1111111101011101 : reciprocal = 1111111111111010;
        16'b1111111101011100 : reciprocal = 1111111111111010;
        16'b1111111101011011 : reciprocal = 1111111111111010;
        16'b1111111101011010 : reciprocal = 1111111111111010;
        16'b1111111101011001 : reciprocal = 1111111111111010;
        16'b1111111101011000 : reciprocal = 1111111111111010;
        16'b1111111101010111 : reciprocal = 1111111111111010;
        16'b1111111101010110 : reciprocal = 1111111111111010;
        16'b1111111101010101 : reciprocal = 1111111111111010;
        16'b1111111101010100 : reciprocal = 1111111111111010;
        16'b1111111101010011 : reciprocal = 1111111111111010;
        16'b1111111101010010 : reciprocal = 1111111111111010;
        16'b1111111101010001 : reciprocal = 1111111111111010;
        16'b1111111101010000 : reciprocal = 1111111111111010;
        16'b1111111101001111 : reciprocal = 1111111111111010;
        16'b1111111101001110 : reciprocal = 1111111111111010;
        16'b1111111101001101 : reciprocal = 1111111111111010;
        16'b1111111101001100 : reciprocal = 1111111111111010;
        16'b1111111101001011 : reciprocal = 1111111111111010;
        16'b1111111101001010 : reciprocal = 1111111111111010;
        16'b1111111101001001 : reciprocal = 1111111111111010;
        16'b1111111101001000 : reciprocal = 1111111111111010;
        16'b1111111101000111 : reciprocal = 1111111111111010;
        16'b1111111101000110 : reciprocal = 1111111111111010;
        16'b1111111101000101 : reciprocal = 1111111111111011;
        16'b1111111101000100 : reciprocal = 1111111111111011;
        16'b1111111101000011 : reciprocal = 1111111111111011;
        16'b1111111101000010 : reciprocal = 1111111111111011;
        16'b1111111101000001 : reciprocal = 1111111111111011;
        16'b1111111101000000 : reciprocal = 1111111111111011;
        16'b1111111100111111 : reciprocal = 1111111111111011;
        16'b1111111100111110 : reciprocal = 1111111111111011;
        16'b1111111100111101 : reciprocal = 1111111111111011;
        16'b1111111100111100 : reciprocal = 1111111111111011;
        16'b1111111100111011 : reciprocal = 1111111111111011;
        16'b1111111100111010 : reciprocal = 1111111111111011;
        16'b1111111100111001 : reciprocal = 1111111111111011;
        16'b1111111100111000 : reciprocal = 1111111111111011;
        16'b1111111100110111 : reciprocal = 1111111111111011;
        16'b1111111100110110 : reciprocal = 1111111111111011;
        16'b1111111100110101 : reciprocal = 1111111111111011;
        16'b1111111100110100 : reciprocal = 1111111111111011;
        16'b1111111100110011 : reciprocal = 1111111111111011;
        16'b1111111100110010 : reciprocal = 1111111111111011;
        16'b1111111100110001 : reciprocal = 1111111111111011;
        16'b1111111100110000 : reciprocal = 1111111111111011;
        16'b1111111100101111 : reciprocal = 1111111111111011;
        16'b1111111100101110 : reciprocal = 1111111111111011;
        16'b1111111100101101 : reciprocal = 1111111111111011;
        16'b1111111100101100 : reciprocal = 1111111111111011;
        16'b1111111100101011 : reciprocal = 1111111111111011;
        16'b1111111100101010 : reciprocal = 1111111111111011;
        16'b1111111100101001 : reciprocal = 1111111111111011;
        16'b1111111100101000 : reciprocal = 1111111111111011;
        16'b1111111100100111 : reciprocal = 1111111111111011;
        16'b1111111100100110 : reciprocal = 1111111111111011;
        16'b1111111100100101 : reciprocal = 1111111111111011;
        16'b1111111100100100 : reciprocal = 1111111111111011;
        16'b1111111100100011 : reciprocal = 1111111111111011;
        16'b1111111100100010 : reciprocal = 1111111111111011;
        16'b1111111100100001 : reciprocal = 1111111111111011;
        16'b1111111100100000 : reciprocal = 1111111111111011;
        16'b1111111100011111 : reciprocal = 1111111111111011;
        16'b1111111100011110 : reciprocal = 1111111111111011;
        16'b1111111100011101 : reciprocal = 1111111111111011;
        16'b1111111100011100 : reciprocal = 1111111111111100;
        16'b1111111100011011 : reciprocal = 1111111111111100;
        16'b1111111100011010 : reciprocal = 1111111111111100;
        16'b1111111100011001 : reciprocal = 1111111111111100;
        16'b1111111100011000 : reciprocal = 1111111111111100;
        16'b1111111100010111 : reciprocal = 1111111111111100;
        16'b1111111100010110 : reciprocal = 1111111111111100;
        16'b1111111100010101 : reciprocal = 1111111111111100;
        16'b1111111100010100 : reciprocal = 1111111111111100;
        16'b1111111100010011 : reciprocal = 1111111111111100;
        16'b1111111100010010 : reciprocal = 1111111111111100;
        16'b1111111100010001 : reciprocal = 1111111111111100;
        16'b1111111100010000 : reciprocal = 1111111111111100;
        16'b1111111100001111 : reciprocal = 1111111111111100;
        16'b1111111100001110 : reciprocal = 1111111111111100;
        16'b1111111100001101 : reciprocal = 1111111111111100;
        16'b1111111100001100 : reciprocal = 1111111111111100;
        16'b1111111100001011 : reciprocal = 1111111111111100;
        16'b1111111100001010 : reciprocal = 1111111111111100;
        16'b1111111100001001 : reciprocal = 1111111111111100;
        16'b1111111100001000 : reciprocal = 1111111111111100;
        16'b1111111100000111 : reciprocal = 1111111111111100;
        16'b1111111100000110 : reciprocal = 1111111111111100;
        16'b1111111100000101 : reciprocal = 1111111111111100;
        16'b1111111100000100 : reciprocal = 1111111111111100;
        16'b1111111100000011 : reciprocal = 1111111111111100;
        16'b1111111100000010 : reciprocal = 1111111111111100;
        16'b1111111100000001 : reciprocal = 1111111111111100;
        16'b1111111100000000 : reciprocal = 1111111111111100;
        16'b1111111011111111 : reciprocal = 1111111111111100;
        16'b1111111011111110 : reciprocal = 1111111111111100;
        16'b1111111011111101 : reciprocal = 1111111111111100;
        16'b1111111011111100 : reciprocal = 1111111111111100;
        16'b1111111011111011 : reciprocal = 1111111111111100;
        16'b1111111011111010 : reciprocal = 1111111111111100;
        16'b1111111011111001 : reciprocal = 1111111111111100;
        16'b1111111011111000 : reciprocal = 1111111111111100;
        16'b1111111011110111 : reciprocal = 1111111111111100;
        16'b1111111011110110 : reciprocal = 1111111111111100;
        16'b1111111011110101 : reciprocal = 1111111111111100;
        16'b1111111011110100 : reciprocal = 1111111111111100;
        16'b1111111011110011 : reciprocal = 1111111111111100;
        16'b1111111011110010 : reciprocal = 1111111111111100;
        16'b1111111011110001 : reciprocal = 1111111111111100;
        16'b1111111011110000 : reciprocal = 1111111111111100;
        16'b1111111011101111 : reciprocal = 1111111111111100;
        16'b1111111011101110 : reciprocal = 1111111111111100;
        16'b1111111011101101 : reciprocal = 1111111111111100;
        16'b1111111011101100 : reciprocal = 1111111111111100;
        16'b1111111011101011 : reciprocal = 1111111111111100;
        16'b1111111011101010 : reciprocal = 1111111111111100;
        16'b1111111011101001 : reciprocal = 1111111111111100;
        16'b1111111011101000 : reciprocal = 1111111111111100;
        16'b1111111011100111 : reciprocal = 1111111111111100;
        16'b1111111011100110 : reciprocal = 1111111111111100;
        16'b1111111011100101 : reciprocal = 1111111111111100;
        16'b1111111011100100 : reciprocal = 1111111111111100;
        16'b1111111011100011 : reciprocal = 1111111111111100;
        16'b1111111011100010 : reciprocal = 1111111111111100;
        16'b1111111011100001 : reciprocal = 1111111111111100;
        16'b1111111011100000 : reciprocal = 1111111111111100;
        16'b1111111011011111 : reciprocal = 1111111111111100;
        16'b1111111011011110 : reciprocal = 1111111111111100;
        16'b1111111011011101 : reciprocal = 1111111111111100;
        16'b1111111011011100 : reciprocal = 1111111111111100;
        16'b1111111011011011 : reciprocal = 1111111111111101;
        16'b1111111011011010 : reciprocal = 1111111111111101;
        16'b1111111011011001 : reciprocal = 1111111111111101;
        16'b1111111011011000 : reciprocal = 1111111111111101;
        16'b1111111011010111 : reciprocal = 1111111111111101;
        16'b1111111011010110 : reciprocal = 1111111111111101;
        16'b1111111011010101 : reciprocal = 1111111111111101;
        16'b1111111011010100 : reciprocal = 1111111111111101;
        16'b1111111011010011 : reciprocal = 1111111111111101;
        16'b1111111011010010 : reciprocal = 1111111111111101;
        16'b1111111011010001 : reciprocal = 1111111111111101;
        16'b1111111011010000 : reciprocal = 1111111111111101;
        16'b1111111011001111 : reciprocal = 1111111111111101;
        16'b1111111011001110 : reciprocal = 1111111111111101;
        16'b1111111011001101 : reciprocal = 1111111111111101;
        16'b1111111011001100 : reciprocal = 1111111111111101;
        16'b1111111011001011 : reciprocal = 1111111111111101;
        16'b1111111011001010 : reciprocal = 1111111111111101;
        16'b1111111011001001 : reciprocal = 1111111111111101;
        16'b1111111011001000 : reciprocal = 1111111111111101;
        16'b1111111011000111 : reciprocal = 1111111111111101;
        16'b1111111011000110 : reciprocal = 1111111111111101;
        16'b1111111011000101 : reciprocal = 1111111111111101;
        16'b1111111011000100 : reciprocal = 1111111111111101;
        16'b1111111011000011 : reciprocal = 1111111111111101;
        16'b1111111011000010 : reciprocal = 1111111111111101;
        16'b1111111011000001 : reciprocal = 1111111111111101;
        16'b1111111011000000 : reciprocal = 1111111111111101;
        16'b1111111010111111 : reciprocal = 1111111111111101;
        16'b1111111010111110 : reciprocal = 1111111111111101;
        16'b1111111010111101 : reciprocal = 1111111111111101;
        16'b1111111010111100 : reciprocal = 1111111111111101;
        16'b1111111010111011 : reciprocal = 1111111111111101;
        16'b1111111010111010 : reciprocal = 1111111111111101;
        16'b1111111010111001 : reciprocal = 1111111111111101;
        16'b1111111010111000 : reciprocal = 1111111111111101;
        16'b1111111010110111 : reciprocal = 1111111111111101;
        16'b1111111010110110 : reciprocal = 1111111111111101;
        16'b1111111010110101 : reciprocal = 1111111111111101;
        16'b1111111010110100 : reciprocal = 1111111111111101;
        16'b1111111010110011 : reciprocal = 1111111111111101;
        16'b1111111010110010 : reciprocal = 1111111111111101;
        16'b1111111010110001 : reciprocal = 1111111111111101;
        16'b1111111010110000 : reciprocal = 1111111111111101;
        16'b1111111010101111 : reciprocal = 1111111111111101;
        16'b1111111010101110 : reciprocal = 1111111111111101;
        16'b1111111010101101 : reciprocal = 1111111111111101;
        16'b1111111010101100 : reciprocal = 1111111111111101;
        16'b1111111010101011 : reciprocal = 1111111111111101;
        16'b1111111010101010 : reciprocal = 1111111111111101;
        16'b1111111010101001 : reciprocal = 1111111111111101;
        16'b1111111010101000 : reciprocal = 1111111111111101;
        16'b1111111010100111 : reciprocal = 1111111111111101;
        16'b1111111010100110 : reciprocal = 1111111111111101;
        16'b1111111010100101 : reciprocal = 1111111111111101;
        16'b1111111010100100 : reciprocal = 1111111111111101;
        16'b1111111010100011 : reciprocal = 1111111111111101;
        16'b1111111010100010 : reciprocal = 1111111111111101;
        16'b1111111010100001 : reciprocal = 1111111111111101;
        16'b1111111010100000 : reciprocal = 1111111111111101;
        16'b1111111010011111 : reciprocal = 1111111111111101;
        16'b1111111010011110 : reciprocal = 1111111111111101;
        16'b1111111010011101 : reciprocal = 1111111111111101;
        16'b1111111010011100 : reciprocal = 1111111111111101;
        16'b1111111010011011 : reciprocal = 1111111111111101;
        16'b1111111010011010 : reciprocal = 1111111111111101;
        16'b1111111010011001 : reciprocal = 1111111111111101;
        16'b1111111010011000 : reciprocal = 1111111111111101;
        16'b1111111010010111 : reciprocal = 1111111111111101;
        16'b1111111010010110 : reciprocal = 1111111111111101;
        16'b1111111010010101 : reciprocal = 1111111111111101;
        16'b1111111010010100 : reciprocal = 1111111111111101;
        16'b1111111010010011 : reciprocal = 1111111111111101;
        16'b1111111010010010 : reciprocal = 1111111111111101;
        16'b1111111010010001 : reciprocal = 1111111111111101;
        16'b1111111010010000 : reciprocal = 1111111111111101;
        16'b1111111010001111 : reciprocal = 1111111111111101;
        16'b1111111010001110 : reciprocal = 1111111111111101;
        16'b1111111010001101 : reciprocal = 1111111111111101;
        16'b1111111010001100 : reciprocal = 1111111111111101;
        16'b1111111010001011 : reciprocal = 1111111111111101;
        16'b1111111010001010 : reciprocal = 1111111111111101;
        16'b1111111010001001 : reciprocal = 1111111111111101;
        16'b1111111010001000 : reciprocal = 1111111111111101;
        16'b1111111010000111 : reciprocal = 1111111111111101;
        16'b1111111010000110 : reciprocal = 1111111111111101;
        16'b1111111010000101 : reciprocal = 1111111111111101;
        16'b1111111010000100 : reciprocal = 1111111111111101;
        16'b1111111010000011 : reciprocal = 1111111111111101;
        16'b1111111010000010 : reciprocal = 1111111111111101;
        16'b1111111010000001 : reciprocal = 1111111111111101;
        16'b1111111010000000 : reciprocal = 1111111111111101;
        16'b1111111001111111 : reciprocal = 1111111111111101;
        16'b1111111001111110 : reciprocal = 1111111111111101;
        16'b1111111001111101 : reciprocal = 1111111111111101;
        16'b1111111001111100 : reciprocal = 1111111111111101;
        16'b1111111001111011 : reciprocal = 1111111111111101;
        16'b1111111001111010 : reciprocal = 1111111111111101;
        16'b1111111001111001 : reciprocal = 1111111111111101;
        16'b1111111001111000 : reciprocal = 1111111111111101;
        16'b1111111001110111 : reciprocal = 1111111111111101;
        16'b1111111001110110 : reciprocal = 1111111111111101;
        16'b1111111001110101 : reciprocal = 1111111111111101;
        16'b1111111001110100 : reciprocal = 1111111111111101;
        16'b1111111001110011 : reciprocal = 1111111111111101;
        16'b1111111001110010 : reciprocal = 1111111111111101;
        16'b1111111001110001 : reciprocal = 1111111111111101;
        16'b1111111001110000 : reciprocal = 1111111111111101;
        16'b1111111001101111 : reciprocal = 1111111111111101;
        16'b1111111001101110 : reciprocal = 1111111111111101;
        16'b1111111001101101 : reciprocal = 1111111111111101;
        16'b1111111001101100 : reciprocal = 1111111111111101;
        16'b1111111001101011 : reciprocal = 1111111111111101;
        16'b1111111001101010 : reciprocal = 1111111111111101;
        16'b1111111001101001 : reciprocal = 1111111111111101;
        16'b1111111001101000 : reciprocal = 1111111111111101;
        16'b1111111001100111 : reciprocal = 1111111111111101;
        16'b1111111001100110 : reciprocal = 1111111111111110;
        16'b1111111001100101 : reciprocal = 1111111111111110;
        16'b1111111001100100 : reciprocal = 1111111111111110;
        16'b1111111001100011 : reciprocal = 1111111111111110;
        16'b1111111001100010 : reciprocal = 1111111111111110;
        16'b1111111001100001 : reciprocal = 1111111111111110;
        16'b1111111001100000 : reciprocal = 1111111111111110;
        16'b1111111001011111 : reciprocal = 1111111111111110;
        16'b1111111001011110 : reciprocal = 1111111111111110;
        16'b1111111001011101 : reciprocal = 1111111111111110;
        16'b1111111001011100 : reciprocal = 1111111111111110;
        16'b1111111001011011 : reciprocal = 1111111111111110;
        16'b1111111001011010 : reciprocal = 1111111111111110;
        16'b1111111001011001 : reciprocal = 1111111111111110;
        16'b1111111001011000 : reciprocal = 1111111111111110;
        16'b1111111001010111 : reciprocal = 1111111111111110;
        16'b1111111001010110 : reciprocal = 1111111111111110;
        16'b1111111001010101 : reciprocal = 1111111111111110;
        16'b1111111001010100 : reciprocal = 1111111111111110;
        16'b1111111001010011 : reciprocal = 1111111111111110;
        16'b1111111001010010 : reciprocal = 1111111111111110;
        16'b1111111001010001 : reciprocal = 1111111111111110;
        16'b1111111001010000 : reciprocal = 1111111111111110;
        16'b1111111001001111 : reciprocal = 1111111111111110;
        16'b1111111001001110 : reciprocal = 1111111111111110;
        16'b1111111001001101 : reciprocal = 1111111111111110;
        16'b1111111001001100 : reciprocal = 1111111111111110;
        16'b1111111001001011 : reciprocal = 1111111111111110;
        16'b1111111001001010 : reciprocal = 1111111111111110;
        16'b1111111001001001 : reciprocal = 1111111111111110;
        16'b1111111001001000 : reciprocal = 1111111111111110;
        16'b1111111001000111 : reciprocal = 1111111111111110;
        16'b1111111001000110 : reciprocal = 1111111111111110;
        16'b1111111001000101 : reciprocal = 1111111111111110;
        16'b1111111001000100 : reciprocal = 1111111111111110;
        16'b1111111001000011 : reciprocal = 1111111111111110;
        16'b1111111001000010 : reciprocal = 1111111111111110;
        16'b1111111001000001 : reciprocal = 1111111111111110;
        16'b1111111001000000 : reciprocal = 1111111111111110;
        16'b1111111000111111 : reciprocal = 1111111111111110;
        16'b1111111000111110 : reciprocal = 1111111111111110;
        16'b1111111000111101 : reciprocal = 1111111111111110;
        16'b1111111000111100 : reciprocal = 1111111111111110;
        16'b1111111000111011 : reciprocal = 1111111111111110;
        16'b1111111000111010 : reciprocal = 1111111111111110;
        16'b1111111000111001 : reciprocal = 1111111111111110;
        16'b1111111000111000 : reciprocal = 1111111111111110;
        16'b1111111000110111 : reciprocal = 1111111111111110;
        16'b1111111000110110 : reciprocal = 1111111111111110;
        16'b1111111000110101 : reciprocal = 1111111111111110;
        16'b1111111000110100 : reciprocal = 1111111111111110;
        16'b1111111000110011 : reciprocal = 1111111111111110;
        16'b1111111000110010 : reciprocal = 1111111111111110;
        16'b1111111000110001 : reciprocal = 1111111111111110;
        16'b1111111000110000 : reciprocal = 1111111111111110;
        16'b1111111000101111 : reciprocal = 1111111111111110;
        16'b1111111000101110 : reciprocal = 1111111111111110;
        16'b1111111000101101 : reciprocal = 1111111111111110;
        16'b1111111000101100 : reciprocal = 1111111111111110;
        16'b1111111000101011 : reciprocal = 1111111111111110;
        16'b1111111000101010 : reciprocal = 1111111111111110;
        16'b1111111000101001 : reciprocal = 1111111111111110;
        16'b1111111000101000 : reciprocal = 1111111111111110;
        16'b1111111000100111 : reciprocal = 1111111111111110;
        16'b1111111000100110 : reciprocal = 1111111111111110;
        16'b1111111000100101 : reciprocal = 1111111111111110;
        16'b1111111000100100 : reciprocal = 1111111111111110;
        16'b1111111000100011 : reciprocal = 1111111111111110;
        16'b1111111000100010 : reciprocal = 1111111111111110;
        16'b1111111000100001 : reciprocal = 1111111111111110;
        16'b1111111000100000 : reciprocal = 1111111111111110;
        16'b1111111000011111 : reciprocal = 1111111111111110;
        16'b1111111000011110 : reciprocal = 1111111111111110;
        16'b1111111000011101 : reciprocal = 1111111111111110;
        16'b1111111000011100 : reciprocal = 1111111111111110;
        16'b1111111000011011 : reciprocal = 1111111111111110;
        16'b1111111000011010 : reciprocal = 1111111111111110;
        16'b1111111000011001 : reciprocal = 1111111111111110;
        16'b1111111000011000 : reciprocal = 1111111111111110;
        16'b1111111000010111 : reciprocal = 1111111111111110;
        16'b1111111000010110 : reciprocal = 1111111111111110;
        16'b1111111000010101 : reciprocal = 1111111111111110;
        16'b1111111000010100 : reciprocal = 1111111111111110;
        16'b1111111000010011 : reciprocal = 1111111111111110;
        16'b1111111000010010 : reciprocal = 1111111111111110;
        16'b1111111000010001 : reciprocal = 1111111111111110;
        16'b1111111000010000 : reciprocal = 1111111111111110;
        16'b1111111000001111 : reciprocal = 1111111111111110;
        16'b1111111000001110 : reciprocal = 1111111111111110;
        16'b1111111000001101 : reciprocal = 1111111111111110;
        16'b1111111000001100 : reciprocal = 1111111111111110;
        16'b1111111000001011 : reciprocal = 1111111111111110;
        16'b1111111000001010 : reciprocal = 1111111111111110;
        16'b1111111000001001 : reciprocal = 1111111111111110;
        16'b1111111000001000 : reciprocal = 1111111111111110;
        16'b1111111000000111 : reciprocal = 1111111111111110;
        16'b1111111000000110 : reciprocal = 1111111111111110;
        16'b1111111000000101 : reciprocal = 1111111111111110;
        16'b1111111000000100 : reciprocal = 1111111111111110;
        16'b1111111000000011 : reciprocal = 1111111111111110;
        16'b1111111000000010 : reciprocal = 1111111111111110;
        16'b1111111000000001 : reciprocal = 1111111111111110;
        16'b1111111000000000 : reciprocal = 1111111111111110;
        16'b1111110111111111 : reciprocal = 1111111111111110;
        16'b1111110111111110 : reciprocal = 1111111111111110;
        16'b1111110111111101 : reciprocal = 1111111111111110;
        16'b1111110111111100 : reciprocal = 1111111111111110;
        16'b1111110111111011 : reciprocal = 1111111111111110;
        16'b1111110111111010 : reciprocal = 1111111111111110;
        16'b1111110111111001 : reciprocal = 1111111111111110;
        16'b1111110111111000 : reciprocal = 1111111111111110;
        16'b1111110111110111 : reciprocal = 1111111111111110;
        16'b1111110111110110 : reciprocal = 1111111111111110;
        16'b1111110111110101 : reciprocal = 1111111111111110;
        16'b1111110111110100 : reciprocal = 1111111111111110;
        16'b1111110111110011 : reciprocal = 1111111111111110;
        16'b1111110111110010 : reciprocal = 1111111111111110;
        16'b1111110111110001 : reciprocal = 1111111111111110;
        16'b1111110111110000 : reciprocal = 1111111111111110;
        16'b1111110111101111 : reciprocal = 1111111111111110;
        16'b1111110111101110 : reciprocal = 1111111111111110;
        16'b1111110111101101 : reciprocal = 1111111111111110;
        16'b1111110111101100 : reciprocal = 1111111111111110;
        16'b1111110111101011 : reciprocal = 1111111111111110;
        16'b1111110111101010 : reciprocal = 1111111111111110;
        16'b1111110111101001 : reciprocal = 1111111111111110;
        16'b1111110111101000 : reciprocal = 1111111111111110;
        16'b1111110111100111 : reciprocal = 1111111111111110;
        16'b1111110111100110 : reciprocal = 1111111111111110;
        16'b1111110111100101 : reciprocal = 1111111111111110;
        16'b1111110111100100 : reciprocal = 1111111111111110;
        16'b1111110111100011 : reciprocal = 1111111111111110;
        16'b1111110111100010 : reciprocal = 1111111111111110;
        16'b1111110111100001 : reciprocal = 1111111111111110;
        16'b1111110111100000 : reciprocal = 1111111111111110;
        16'b1111110111011111 : reciprocal = 1111111111111110;
        16'b1111110111011110 : reciprocal = 1111111111111110;
        16'b1111110111011101 : reciprocal = 1111111111111110;
        16'b1111110111011100 : reciprocal = 1111111111111110;
        16'b1111110111011011 : reciprocal = 1111111111111110;
        16'b1111110111011010 : reciprocal = 1111111111111110;
        16'b1111110111011001 : reciprocal = 1111111111111110;
        16'b1111110111011000 : reciprocal = 1111111111111110;
        16'b1111110111010111 : reciprocal = 1111111111111110;
        16'b1111110111010110 : reciprocal = 1111111111111110;
        16'b1111110111010101 : reciprocal = 1111111111111110;
        16'b1111110111010100 : reciprocal = 1111111111111110;
        16'b1111110111010011 : reciprocal = 1111111111111110;
        16'b1111110111010010 : reciprocal = 1111111111111110;
        16'b1111110111010001 : reciprocal = 1111111111111110;
        16'b1111110111010000 : reciprocal = 1111111111111110;
        16'b1111110111001111 : reciprocal = 1111111111111110;
        16'b1111110111001110 : reciprocal = 1111111111111110;
        16'b1111110111001101 : reciprocal = 1111111111111110;
        16'b1111110111001100 : reciprocal = 1111111111111110;
        16'b1111110111001011 : reciprocal = 1111111111111110;
        16'b1111110111001010 : reciprocal = 1111111111111110;
        16'b1111110111001001 : reciprocal = 1111111111111110;
        16'b1111110111001000 : reciprocal = 1111111111111110;
        16'b1111110111000111 : reciprocal = 1111111111111110;
        16'b1111110111000110 : reciprocal = 1111111111111110;
        16'b1111110111000101 : reciprocal = 1111111111111110;
        16'b1111110111000100 : reciprocal = 1111111111111110;
        16'b1111110111000011 : reciprocal = 1111111111111110;
        16'b1111110111000010 : reciprocal = 1111111111111110;
        16'b1111110111000001 : reciprocal = 1111111111111110;
        16'b1111110111000000 : reciprocal = 1111111111111110;
        16'b1111110110111111 : reciprocal = 1111111111111110;
        16'b1111110110111110 : reciprocal = 1111111111111110;
        16'b1111110110111101 : reciprocal = 1111111111111110;
        16'b1111110110111100 : reciprocal = 1111111111111110;
        16'b1111110110111011 : reciprocal = 1111111111111110;
        16'b1111110110111010 : reciprocal = 1111111111111110;
        16'b1111110110111001 : reciprocal = 1111111111111110;
        16'b1111110110111000 : reciprocal = 1111111111111110;
        16'b1111110110110111 : reciprocal = 1111111111111110;
        16'b1111110110110110 : reciprocal = 1111111111111110;
        16'b1111110110110101 : reciprocal = 1111111111111110;
        16'b1111110110110100 : reciprocal = 1111111111111110;
        16'b1111110110110011 : reciprocal = 1111111111111110;
        16'b1111110110110010 : reciprocal = 1111111111111110;
        16'b1111110110110001 : reciprocal = 1111111111111110;
        16'b1111110110110000 : reciprocal = 1111111111111110;
        16'b1111110110101111 : reciprocal = 1111111111111110;
        16'b1111110110101110 : reciprocal = 1111111111111110;
        16'b1111110110101101 : reciprocal = 1111111111111110;
        16'b1111110110101100 : reciprocal = 1111111111111110;
        16'b1111110110101011 : reciprocal = 1111111111111110;
        16'b1111110110101010 : reciprocal = 1111111111111110;
        16'b1111110110101001 : reciprocal = 1111111111111110;
        16'b1111110110101000 : reciprocal = 1111111111111110;
        16'b1111110110100111 : reciprocal = 1111111111111110;
        16'b1111110110100110 : reciprocal = 1111111111111110;
        16'b1111110110100101 : reciprocal = 1111111111111110;
        16'b1111110110100100 : reciprocal = 1111111111111110;
        16'b1111110110100011 : reciprocal = 1111111111111110;
        16'b1111110110100010 : reciprocal = 1111111111111110;
        16'b1111110110100001 : reciprocal = 1111111111111110;
        16'b1111110110100000 : reciprocal = 1111111111111110;
        16'b1111110110011111 : reciprocal = 1111111111111110;
        16'b1111110110011110 : reciprocal = 1111111111111110;
        16'b1111110110011101 : reciprocal = 1111111111111110;
        16'b1111110110011100 : reciprocal = 1111111111111110;
        16'b1111110110011011 : reciprocal = 1111111111111110;
        16'b1111110110011010 : reciprocal = 1111111111111110;
        16'b1111110110011001 : reciprocal = 1111111111111110;
        16'b1111110110011000 : reciprocal = 1111111111111110;
        16'b1111110110010111 : reciprocal = 1111111111111110;
        16'b1111110110010110 : reciprocal = 1111111111111110;
        16'b1111110110010101 : reciprocal = 1111111111111110;
        16'b1111110110010100 : reciprocal = 1111111111111110;
        16'b1111110110010011 : reciprocal = 1111111111111110;
        16'b1111110110010010 : reciprocal = 1111111111111110;
        16'b1111110110010001 : reciprocal = 1111111111111110;
        16'b1111110110010000 : reciprocal = 1111111111111110;
        16'b1111110110001111 : reciprocal = 1111111111111110;
        16'b1111110110001110 : reciprocal = 1111111111111110;
        16'b1111110110001101 : reciprocal = 1111111111111110;
        16'b1111110110001100 : reciprocal = 1111111111111110;
        16'b1111110110001011 : reciprocal = 1111111111111110;
        16'b1111110110001010 : reciprocal = 1111111111111110;
        16'b1111110110001001 : reciprocal = 1111111111111110;
        16'b1111110110001000 : reciprocal = 1111111111111110;
        16'b1111110110000111 : reciprocal = 1111111111111110;
        16'b1111110110000110 : reciprocal = 1111111111111110;
        16'b1111110110000101 : reciprocal = 1111111111111110;
        16'b1111110110000100 : reciprocal = 1111111111111110;
        16'b1111110110000011 : reciprocal = 1111111111111110;
        16'b1111110110000010 : reciprocal = 1111111111111110;
        16'b1111110110000001 : reciprocal = 1111111111111110;
        16'b1111110110000000 : reciprocal = 1111111111111110;
        16'b1111110101111111 : reciprocal = 1111111111111110;
        16'b1111110101111110 : reciprocal = 1111111111111110;
        16'b1111110101111101 : reciprocal = 1111111111111110;
        16'b1111110101111100 : reciprocal = 1111111111111110;
        16'b1111110101111011 : reciprocal = 1111111111111110;
        16'b1111110101111010 : reciprocal = 1111111111111110;
        16'b1111110101111001 : reciprocal = 1111111111111110;
        16'b1111110101111000 : reciprocal = 1111111111111110;
        16'b1111110101110111 : reciprocal = 1111111111111110;
        16'b1111110101110110 : reciprocal = 1111111111111110;
        16'b1111110101110101 : reciprocal = 1111111111111110;
        16'b1111110101110100 : reciprocal = 1111111111111110;
        16'b1111110101110011 : reciprocal = 1111111111111110;
        16'b1111110101110010 : reciprocal = 1111111111111110;
        16'b1111110101110001 : reciprocal = 1111111111111110;
        16'b1111110101110000 : reciprocal = 1111111111111110;
        16'b1111110101101111 : reciprocal = 1111111111111110;
        16'b1111110101101110 : reciprocal = 1111111111111110;
        16'b1111110101101101 : reciprocal = 1111111111111110;
        16'b1111110101101100 : reciprocal = 1111111111111110;
        16'b1111110101101011 : reciprocal = 1111111111111110;
        16'b1111110101101010 : reciprocal = 1111111111111110;
        16'b1111110101101001 : reciprocal = 1111111111111110;
        16'b1111110101101000 : reciprocal = 1111111111111110;
        16'b1111110101100111 : reciprocal = 1111111111111110;
        16'b1111110101100110 : reciprocal = 1111111111111110;
        16'b1111110101100101 : reciprocal = 1111111111111110;
        16'b1111110101100100 : reciprocal = 1111111111111110;
        16'b1111110101100011 : reciprocal = 1111111111111110;
        16'b1111110101100010 : reciprocal = 1111111111111110;
        16'b1111110101100001 : reciprocal = 1111111111111110;
        16'b1111110101100000 : reciprocal = 1111111111111110;
        16'b1111110101011111 : reciprocal = 1111111111111110;
        16'b1111110101011110 : reciprocal = 1111111111111110;
        16'b1111110101011101 : reciprocal = 1111111111111110;
        16'b1111110101011100 : reciprocal = 1111111111111110;
        16'b1111110101011011 : reciprocal = 1111111111111110;
        16'b1111110101011010 : reciprocal = 1111111111111110;
        16'b1111110101011001 : reciprocal = 1111111111111110;
        16'b1111110101011000 : reciprocal = 1111111111111110;
        16'b1111110101010111 : reciprocal = 1111111111111110;
        16'b1111110101010110 : reciprocal = 1111111111111110;
        16'b1111110101010101 : reciprocal = 1111111111111111;
        16'b1111110101010100 : reciprocal = 1111111111111111;
        16'b1111110101010011 : reciprocal = 1111111111111111;
        16'b1111110101010010 : reciprocal = 1111111111111111;
        16'b1111110101010001 : reciprocal = 1111111111111111;
        16'b1111110101010000 : reciprocal = 1111111111111111;
        16'b1111110101001111 : reciprocal = 1111111111111111;
        16'b1111110101001110 : reciprocal = 1111111111111111;
        16'b1111110101001101 : reciprocal = 1111111111111111;
        16'b1111110101001100 : reciprocal = 1111111111111111;
        16'b1111110101001011 : reciprocal = 1111111111111111;
        16'b1111110101001010 : reciprocal = 1111111111111111;
        16'b1111110101001001 : reciprocal = 1111111111111111;
        16'b1111110101001000 : reciprocal = 1111111111111111;
        16'b1111110101000111 : reciprocal = 1111111111111111;
        16'b1111110101000110 : reciprocal = 1111111111111111;
        16'b1111110101000101 : reciprocal = 1111111111111111;
        16'b1111110101000100 : reciprocal = 1111111111111111;
        16'b1111110101000011 : reciprocal = 1111111111111111;
        16'b1111110101000010 : reciprocal = 1111111111111111;
        16'b1111110101000001 : reciprocal = 1111111111111111;
        16'b1111110101000000 : reciprocal = 1111111111111111;
        16'b1111110100111111 : reciprocal = 1111111111111111;
        16'b1111110100111110 : reciprocal = 1111111111111111;
        16'b1111110100111101 : reciprocal = 1111111111111111;
        16'b1111110100111100 : reciprocal = 1111111111111111;
        16'b1111110100111011 : reciprocal = 1111111111111111;
        16'b1111110100111010 : reciprocal = 1111111111111111;
        16'b1111110100111001 : reciprocal = 1111111111111111;
        16'b1111110100111000 : reciprocal = 1111111111111111;
        16'b1111110100110111 : reciprocal = 1111111111111111;
        16'b1111110100110110 : reciprocal = 1111111111111111;
        16'b1111110100110101 : reciprocal = 1111111111111111;
        16'b1111110100110100 : reciprocal = 1111111111111111;
        16'b1111110100110011 : reciprocal = 1111111111111111;
        16'b1111110100110010 : reciprocal = 1111111111111111;
        16'b1111110100110001 : reciprocal = 1111111111111111;
        16'b1111110100110000 : reciprocal = 1111111111111111;
        16'b1111110100101111 : reciprocal = 1111111111111111;
        16'b1111110100101110 : reciprocal = 1111111111111111;
        16'b1111110100101101 : reciprocal = 1111111111111111;
        16'b1111110100101100 : reciprocal = 1111111111111111;
        16'b1111110100101011 : reciprocal = 1111111111111111;
        16'b1111110100101010 : reciprocal = 1111111111111111;
        16'b1111110100101001 : reciprocal = 1111111111111111;
        16'b1111110100101000 : reciprocal = 1111111111111111;
        16'b1111110100100111 : reciprocal = 1111111111111111;
        16'b1111110100100110 : reciprocal = 1111111111111111;
        16'b1111110100100101 : reciprocal = 1111111111111111;
        16'b1111110100100100 : reciprocal = 1111111111111111;
        16'b1111110100100011 : reciprocal = 1111111111111111;
        16'b1111110100100010 : reciprocal = 1111111111111111;
        16'b1111110100100001 : reciprocal = 1111111111111111;
        16'b1111110100100000 : reciprocal = 1111111111111111;
        16'b1111110100011111 : reciprocal = 1111111111111111;
        16'b1111110100011110 : reciprocal = 1111111111111111;
        16'b1111110100011101 : reciprocal = 1111111111111111;
        16'b1111110100011100 : reciprocal = 1111111111111111;
        16'b1111110100011011 : reciprocal = 1111111111111111;
        16'b1111110100011010 : reciprocal = 1111111111111111;
        16'b1111110100011001 : reciprocal = 1111111111111111;
        16'b1111110100011000 : reciprocal = 1111111111111111;
        16'b1111110100010111 : reciprocal = 1111111111111111;
        16'b1111110100010110 : reciprocal = 1111111111111111;
        16'b1111110100010101 : reciprocal = 1111111111111111;
        16'b1111110100010100 : reciprocal = 1111111111111111;
        16'b1111110100010011 : reciprocal = 1111111111111111;
        16'b1111110100010010 : reciprocal = 1111111111111111;
        16'b1111110100010001 : reciprocal = 1111111111111111;
        16'b1111110100010000 : reciprocal = 1111111111111111;
        16'b1111110100001111 : reciprocal = 1111111111111111;
        16'b1111110100001110 : reciprocal = 1111111111111111;
        16'b1111110100001101 : reciprocal = 1111111111111111;
        16'b1111110100001100 : reciprocal = 1111111111111111;
        16'b1111110100001011 : reciprocal = 1111111111111111;
        16'b1111110100001010 : reciprocal = 1111111111111111;
        16'b1111110100001001 : reciprocal = 1111111111111111;
        16'b1111110100001000 : reciprocal = 1111111111111111;
        16'b1111110100000111 : reciprocal = 1111111111111111;
        16'b1111110100000110 : reciprocal = 1111111111111111;
        16'b1111110100000101 : reciprocal = 1111111111111111;
        16'b1111110100000100 : reciprocal = 1111111111111111;
        16'b1111110100000011 : reciprocal = 1111111111111111;
        16'b1111110100000010 : reciprocal = 1111111111111111;
        16'b1111110100000001 : reciprocal = 1111111111111111;
        16'b1111110100000000 : reciprocal = 1111111111111111;
        16'b1111110011111111 : reciprocal = 1111111111111111;
        16'b1111110011111110 : reciprocal = 1111111111111111;
        16'b1111110011111101 : reciprocal = 1111111111111111;
        16'b1111110011111100 : reciprocal = 1111111111111111;
        16'b1111110011111011 : reciprocal = 1111111111111111;
        16'b1111110011111010 : reciprocal = 1111111111111111;
        16'b1111110011111001 : reciprocal = 1111111111111111;
        16'b1111110011111000 : reciprocal = 1111111111111111;
        16'b1111110011110111 : reciprocal = 1111111111111111;
        16'b1111110011110110 : reciprocal = 1111111111111111;
        16'b1111110011110101 : reciprocal = 1111111111111111;
        16'b1111110011110100 : reciprocal = 1111111111111111;
        16'b1111110011110011 : reciprocal = 1111111111111111;
        16'b1111110011110010 : reciprocal = 1111111111111111;
        16'b1111110011110001 : reciprocal = 1111111111111111;
        16'b1111110011110000 : reciprocal = 1111111111111111;
        16'b1111110011101111 : reciprocal = 1111111111111111;
        16'b1111110011101110 : reciprocal = 1111111111111111;
        16'b1111110011101101 : reciprocal = 1111111111111111;
        16'b1111110011101100 : reciprocal = 1111111111111111;
        16'b1111110011101011 : reciprocal = 1111111111111111;
        16'b1111110011101010 : reciprocal = 1111111111111111;
        16'b1111110011101001 : reciprocal = 1111111111111111;
        16'b1111110011101000 : reciprocal = 1111111111111111;
        16'b1111110011100111 : reciprocal = 1111111111111111;
        16'b1111110011100110 : reciprocal = 1111111111111111;
        16'b1111110011100101 : reciprocal = 1111111111111111;
        16'b1111110011100100 : reciprocal = 1111111111111111;
        16'b1111110011100011 : reciprocal = 1111111111111111;
        16'b1111110011100010 : reciprocal = 1111111111111111;
        16'b1111110011100001 : reciprocal = 1111111111111111;
        16'b1111110011100000 : reciprocal = 1111111111111111;
        16'b1111110011011111 : reciprocal = 1111111111111111;
        16'b1111110011011110 : reciprocal = 1111111111111111;
        16'b1111110011011101 : reciprocal = 1111111111111111;
        16'b1111110011011100 : reciprocal = 1111111111111111;
        16'b1111110011011011 : reciprocal = 1111111111111111;
        16'b1111110011011010 : reciprocal = 1111111111111111;
        16'b1111110011011001 : reciprocal = 1111111111111111;
        16'b1111110011011000 : reciprocal = 1111111111111111;
        16'b1111110011010111 : reciprocal = 1111111111111111;
        16'b1111110011010110 : reciprocal = 1111111111111111;
        16'b1111110011010101 : reciprocal = 1111111111111111;
        16'b1111110011010100 : reciprocal = 1111111111111111;
        16'b1111110011010011 : reciprocal = 1111111111111111;
        16'b1111110011010010 : reciprocal = 1111111111111111;
        16'b1111110011010001 : reciprocal = 1111111111111111;
        16'b1111110011010000 : reciprocal = 1111111111111111;
        16'b1111110011001111 : reciprocal = 1111111111111111;
        16'b1111110011001110 : reciprocal = 1111111111111111;
        16'b1111110011001101 : reciprocal = 1111111111111111;
        16'b1111110011001100 : reciprocal = 1111111111111111;
        16'b1111110011001011 : reciprocal = 1111111111111111;
        16'b1111110011001010 : reciprocal = 1111111111111111;
        16'b1111110011001001 : reciprocal = 1111111111111111;
        16'b1111110011001000 : reciprocal = 1111111111111111;
        16'b1111110011000111 : reciprocal = 1111111111111111;
        16'b1111110011000110 : reciprocal = 1111111111111111;
        16'b1111110011000101 : reciprocal = 1111111111111111;
        16'b1111110011000100 : reciprocal = 1111111111111111;
        16'b1111110011000011 : reciprocal = 1111111111111111;
        16'b1111110011000010 : reciprocal = 1111111111111111;
        16'b1111110011000001 : reciprocal = 1111111111111111;
        16'b1111110011000000 : reciprocal = 1111111111111111;
        16'b1111110010111111 : reciprocal = 1111111111111111;
        16'b1111110010111110 : reciprocal = 1111111111111111;
        16'b1111110010111101 : reciprocal = 1111111111111111;
        16'b1111110010111100 : reciprocal = 1111111111111111;
        16'b1111110010111011 : reciprocal = 1111111111111111;
        16'b1111110010111010 : reciprocal = 1111111111111111;
        16'b1111110010111001 : reciprocal = 1111111111111111;
        16'b1111110010111000 : reciprocal = 1111111111111111;
        16'b1111110010110111 : reciprocal = 1111111111111111;
        16'b1111110010110110 : reciprocal = 1111111111111111;
        16'b1111110010110101 : reciprocal = 1111111111111111;
        16'b1111110010110100 : reciprocal = 1111111111111111;
        16'b1111110010110011 : reciprocal = 1111111111111111;
        16'b1111110010110010 : reciprocal = 1111111111111111;
        16'b1111110010110001 : reciprocal = 1111111111111111;
        16'b1111110010110000 : reciprocal = 1111111111111111;
        16'b1111110010101111 : reciprocal = 1111111111111111;
        16'b1111110010101110 : reciprocal = 1111111111111111;
        16'b1111110010101101 : reciprocal = 1111111111111111;
        16'b1111110010101100 : reciprocal = 1111111111111111;
        16'b1111110010101011 : reciprocal = 1111111111111111;
        16'b1111110010101010 : reciprocal = 1111111111111111;
        16'b1111110010101001 : reciprocal = 1111111111111111;
        16'b1111110010101000 : reciprocal = 1111111111111111;
        16'b1111110010100111 : reciprocal = 1111111111111111;
        16'b1111110010100110 : reciprocal = 1111111111111111;
        16'b1111110010100101 : reciprocal = 1111111111111111;
        16'b1111110010100100 : reciprocal = 1111111111111111;
        16'b1111110010100011 : reciprocal = 1111111111111111;
        16'b1111110010100010 : reciprocal = 1111111111111111;
        16'b1111110010100001 : reciprocal = 1111111111111111;
        16'b1111110010100000 : reciprocal = 1111111111111111;
        16'b1111110010011111 : reciprocal = 1111111111111111;
        16'b1111110010011110 : reciprocal = 1111111111111111;
        16'b1111110010011101 : reciprocal = 1111111111111111;
        16'b1111110010011100 : reciprocal = 1111111111111111;
        16'b1111110010011011 : reciprocal = 1111111111111111;
        16'b1111110010011010 : reciprocal = 1111111111111111;
        16'b1111110010011001 : reciprocal = 1111111111111111;
        16'b1111110010011000 : reciprocal = 1111111111111111;
        16'b1111110010010111 : reciprocal = 1111111111111111;
        16'b1111110010010110 : reciprocal = 1111111111111111;
        16'b1111110010010101 : reciprocal = 1111111111111111;
        16'b1111110010010100 : reciprocal = 1111111111111111;
        16'b1111110010010011 : reciprocal = 1111111111111111;
        16'b1111110010010010 : reciprocal = 1111111111111111;
        16'b1111110010010001 : reciprocal = 1111111111111111;
        16'b1111110010010000 : reciprocal = 1111111111111111;
        16'b1111110010001111 : reciprocal = 1111111111111111;
        16'b1111110010001110 : reciprocal = 1111111111111111;
        16'b1111110010001101 : reciprocal = 1111111111111111;
        16'b1111110010001100 : reciprocal = 1111111111111111;
        16'b1111110010001011 : reciprocal = 1111111111111111;
        16'b1111110010001010 : reciprocal = 1111111111111111;
        16'b1111110010001001 : reciprocal = 1111111111111111;
        16'b1111110010001000 : reciprocal = 1111111111111111;
        16'b1111110010000111 : reciprocal = 1111111111111111;
        16'b1111110010000110 : reciprocal = 1111111111111111;
        16'b1111110010000101 : reciprocal = 1111111111111111;
        16'b1111110010000100 : reciprocal = 1111111111111111;
        16'b1111110010000011 : reciprocal = 1111111111111111;
        16'b1111110010000010 : reciprocal = 1111111111111111;
        16'b1111110010000001 : reciprocal = 1111111111111111;
        16'b1111110010000000 : reciprocal = 1111111111111111;
        16'b1111110001111111 : reciprocal = 1111111111111111;
        16'b1111110001111110 : reciprocal = 1111111111111111;
        16'b1111110001111101 : reciprocal = 1111111111111111;
        16'b1111110001111100 : reciprocal = 1111111111111111;
        16'b1111110001111011 : reciprocal = 1111111111111111;
        16'b1111110001111010 : reciprocal = 1111111111111111;
        16'b1111110001111001 : reciprocal = 1111111111111111;
        16'b1111110001111000 : reciprocal = 1111111111111111;
        16'b1111110001110111 : reciprocal = 1111111111111111;
        16'b1111110001110110 : reciprocal = 1111111111111111;
        16'b1111110001110101 : reciprocal = 1111111111111111;
        16'b1111110001110100 : reciprocal = 1111111111111111;
        16'b1111110001110011 : reciprocal = 1111111111111111;
        16'b1111110001110010 : reciprocal = 1111111111111111;
        16'b1111110001110001 : reciprocal = 1111111111111111;
        16'b1111110001110000 : reciprocal = 1111111111111111;
        16'b1111110001101111 : reciprocal = 1111111111111111;
        16'b1111110001101110 : reciprocal = 1111111111111111;
        16'b1111110001101101 : reciprocal = 1111111111111111;
        16'b1111110001101100 : reciprocal = 1111111111111111;
        16'b1111110001101011 : reciprocal = 1111111111111111;
        16'b1111110001101010 : reciprocal = 1111111111111111;
        16'b1111110001101001 : reciprocal = 1111111111111111;
        16'b1111110001101000 : reciprocal = 1111111111111111;
        16'b1111110001100111 : reciprocal = 1111111111111111;
        16'b1111110001100110 : reciprocal = 1111111111111111;
        16'b1111110001100101 : reciprocal = 1111111111111111;
        16'b1111110001100100 : reciprocal = 1111111111111111;
        16'b1111110001100011 : reciprocal = 1111111111111111;
        16'b1111110001100010 : reciprocal = 1111111111111111;
        16'b1111110001100001 : reciprocal = 1111111111111111;
        16'b1111110001100000 : reciprocal = 1111111111111111;
        16'b1111110001011111 : reciprocal = 1111111111111111;
        16'b1111110001011110 : reciprocal = 1111111111111111;
        16'b1111110001011101 : reciprocal = 1111111111111111;
        16'b1111110001011100 : reciprocal = 1111111111111111;
        16'b1111110001011011 : reciprocal = 1111111111111111;
        16'b1111110001011010 : reciprocal = 1111111111111111;
        16'b1111110001011001 : reciprocal = 1111111111111111;
        16'b1111110001011000 : reciprocal = 1111111111111111;
        16'b1111110001010111 : reciprocal = 1111111111111111;
        16'b1111110001010110 : reciprocal = 1111111111111111;
        16'b1111110001010101 : reciprocal = 1111111111111111;
        16'b1111110001010100 : reciprocal = 1111111111111111;
        16'b1111110001010011 : reciprocal = 1111111111111111;
        16'b1111110001010010 : reciprocal = 1111111111111111;
        16'b1111110001010001 : reciprocal = 1111111111111111;
        16'b1111110001010000 : reciprocal = 1111111111111111;
        16'b1111110001001111 : reciprocal = 1111111111111111;
        16'b1111110001001110 : reciprocal = 1111111111111111;
        16'b1111110001001101 : reciprocal = 1111111111111111;
        16'b1111110001001100 : reciprocal = 1111111111111111;
        16'b1111110001001011 : reciprocal = 1111111111111111;
        16'b1111110001001010 : reciprocal = 1111111111111111;
        16'b1111110001001001 : reciprocal = 1111111111111111;
        16'b1111110001001000 : reciprocal = 1111111111111111;
        16'b1111110001000111 : reciprocal = 1111111111111111;
        16'b1111110001000110 : reciprocal = 1111111111111111;
        16'b1111110001000101 : reciprocal = 1111111111111111;
        16'b1111110001000100 : reciprocal = 1111111111111111;
        16'b1111110001000011 : reciprocal = 1111111111111111;
        16'b1111110001000010 : reciprocal = 1111111111111111;
        16'b1111110001000001 : reciprocal = 1111111111111111;
        16'b1111110001000000 : reciprocal = 1111111111111111;
        16'b1111110000111111 : reciprocal = 1111111111111111;
        16'b1111110000111110 : reciprocal = 1111111111111111;
        16'b1111110000111101 : reciprocal = 1111111111111111;
        16'b1111110000111100 : reciprocal = 1111111111111111;
        16'b1111110000111011 : reciprocal = 1111111111111111;
        16'b1111110000111010 : reciprocal = 1111111111111111;
        16'b1111110000111001 : reciprocal = 1111111111111111;
        16'b1111110000111000 : reciprocal = 1111111111111111;
        16'b1111110000110111 : reciprocal = 1111111111111111;
        16'b1111110000110110 : reciprocal = 1111111111111111;
        16'b1111110000110101 : reciprocal = 1111111111111111;
        16'b1111110000110100 : reciprocal = 1111111111111111;
        16'b1111110000110011 : reciprocal = 1111111111111111;
        16'b1111110000110010 : reciprocal = 1111111111111111;
        16'b1111110000110001 : reciprocal = 1111111111111111;
        16'b1111110000110000 : reciprocal = 1111111111111111;
        16'b1111110000101111 : reciprocal = 1111111111111111;
        16'b1111110000101110 : reciprocal = 1111111111111111;
        16'b1111110000101101 : reciprocal = 1111111111111111;
        16'b1111110000101100 : reciprocal = 1111111111111111;
        16'b1111110000101011 : reciprocal = 1111111111111111;
        16'b1111110000101010 : reciprocal = 1111111111111111;
        16'b1111110000101001 : reciprocal = 1111111111111111;
        16'b1111110000101000 : reciprocal = 1111111111111111;
        16'b1111110000100111 : reciprocal = 1111111111111111;
        16'b1111110000100110 : reciprocal = 1111111111111111;
        16'b1111110000100101 : reciprocal = 1111111111111111;
        16'b1111110000100100 : reciprocal = 1111111111111111;
        16'b1111110000100011 : reciprocal = 1111111111111111;
        16'b1111110000100010 : reciprocal = 1111111111111111;
        16'b1111110000100001 : reciprocal = 1111111111111111;
        16'b1111110000100000 : reciprocal = 1111111111111111;
        16'b1111110000011111 : reciprocal = 1111111111111111;
        16'b1111110000011110 : reciprocal = 1111111111111111;
        16'b1111110000011101 : reciprocal = 1111111111111111;
        16'b1111110000011100 : reciprocal = 1111111111111111;
        16'b1111110000011011 : reciprocal = 1111111111111111;
        16'b1111110000011010 : reciprocal = 1111111111111111;
        16'b1111110000011001 : reciprocal = 1111111111111111;
        16'b1111110000011000 : reciprocal = 1111111111111111;
        16'b1111110000010111 : reciprocal = 1111111111111111;
        16'b1111110000010110 : reciprocal = 1111111111111111;
        16'b1111110000010101 : reciprocal = 1111111111111111;
        16'b1111110000010100 : reciprocal = 1111111111111111;
        16'b1111110000010011 : reciprocal = 1111111111111111;
        16'b1111110000010010 : reciprocal = 1111111111111111;
        16'b1111110000010001 : reciprocal = 1111111111111111;
        16'b1111110000010000 : reciprocal = 1111111111111111;
        16'b1111110000001111 : reciprocal = 1111111111111111;
        16'b1111110000001110 : reciprocal = 1111111111111111;
        16'b1111110000001101 : reciprocal = 1111111111111111;
        16'b1111110000001100 : reciprocal = 1111111111111111;
        16'b1111110000001011 : reciprocal = 1111111111111111;
        16'b1111110000001010 : reciprocal = 1111111111111111;
        16'b1111110000001001 : reciprocal = 1111111111111111;
        16'b1111110000001000 : reciprocal = 1111111111111111;
        16'b1111110000000111 : reciprocal = 1111111111111111;
        16'b1111110000000110 : reciprocal = 1111111111111111;
        16'b1111110000000101 : reciprocal = 1111111111111111;
        16'b1111110000000100 : reciprocal = 1111111111111111;
        16'b1111110000000011 : reciprocal = 1111111111111111;
        16'b1111110000000010 : reciprocal = 1111111111111111;
        16'b1111110000000001 : reciprocal = 1111111111111111;
        16'b1111110000000000 : reciprocal = 1111111111111111;
        16'b1111101111111111 : reciprocal = 1111111111111111;
        16'b1111101111111110 : reciprocal = 1111111111111111;
        16'b1111101111111101 : reciprocal = 1111111111111111;
        16'b1111101111111100 : reciprocal = 1111111111111111;
        16'b1111101111111011 : reciprocal = 1111111111111111;
        16'b1111101111111010 : reciprocal = 1111111111111111;
        16'b1111101111111001 : reciprocal = 1111111111111111;
        16'b1111101111111000 : reciprocal = 1111111111111111;
        16'b1111101111110111 : reciprocal = 1111111111111111;
        16'b1111101111110110 : reciprocal = 1111111111111111;
        16'b1111101111110101 : reciprocal = 1111111111111111;
        16'b1111101111110100 : reciprocal = 1111111111111111;
        16'b1111101111110011 : reciprocal = 1111111111111111;
        16'b1111101111110010 : reciprocal = 1111111111111111;
        16'b1111101111110001 : reciprocal = 1111111111111111;
        16'b1111101111110000 : reciprocal = 1111111111111111;
        16'b1111101111101111 : reciprocal = 1111111111111111;
        16'b1111101111101110 : reciprocal = 1111111111111111;
        16'b1111101111101101 : reciprocal = 1111111111111111;
        16'b1111101111101100 : reciprocal = 1111111111111111;
        16'b1111101111101011 : reciprocal = 1111111111111111;
        16'b1111101111101010 : reciprocal = 1111111111111111;
        16'b1111101111101001 : reciprocal = 1111111111111111;
        16'b1111101111101000 : reciprocal = 1111111111111111;
        16'b1111101111100111 : reciprocal = 1111111111111111;
        16'b1111101111100110 : reciprocal = 1111111111111111;
        16'b1111101111100101 : reciprocal = 1111111111111111;
        16'b1111101111100100 : reciprocal = 1111111111111111;
        16'b1111101111100011 : reciprocal = 1111111111111111;
        16'b1111101111100010 : reciprocal = 1111111111111111;
        16'b1111101111100001 : reciprocal = 1111111111111111;
        16'b1111101111100000 : reciprocal = 1111111111111111;
        16'b1111101111011111 : reciprocal = 1111111111111111;
        16'b1111101111011110 : reciprocal = 1111111111111111;
        16'b1111101111011101 : reciprocal = 1111111111111111;
        16'b1111101111011100 : reciprocal = 1111111111111111;
        16'b1111101111011011 : reciprocal = 1111111111111111;
        16'b1111101111011010 : reciprocal = 1111111111111111;
        16'b1111101111011001 : reciprocal = 1111111111111111;
        16'b1111101111011000 : reciprocal = 1111111111111111;
        16'b1111101111010111 : reciprocal = 1111111111111111;
        16'b1111101111010110 : reciprocal = 1111111111111111;
        16'b1111101111010101 : reciprocal = 1111111111111111;
        16'b1111101111010100 : reciprocal = 1111111111111111;
        16'b1111101111010011 : reciprocal = 1111111111111111;
        16'b1111101111010010 : reciprocal = 1111111111111111;
        16'b1111101111010001 : reciprocal = 1111111111111111;
        16'b1111101111010000 : reciprocal = 1111111111111111;
        16'b1111101111001111 : reciprocal = 1111111111111111;
        16'b1111101111001110 : reciprocal = 1111111111111111;
        16'b1111101111001101 : reciprocal = 1111111111111111;
        16'b1111101111001100 : reciprocal = 1111111111111111;
        16'b1111101111001011 : reciprocal = 1111111111111111;
        16'b1111101111001010 : reciprocal = 1111111111111111;
        16'b1111101111001001 : reciprocal = 1111111111111111;
        16'b1111101111001000 : reciprocal = 1111111111111111;
        16'b1111101111000111 : reciprocal = 1111111111111111;
        16'b1111101111000110 : reciprocal = 1111111111111111;
        16'b1111101111000101 : reciprocal = 1111111111111111;
        16'b1111101111000100 : reciprocal = 1111111111111111;
        16'b1111101111000011 : reciprocal = 1111111111111111;
        16'b1111101111000010 : reciprocal = 1111111111111111;
        16'b1111101111000001 : reciprocal = 1111111111111111;
        16'b1111101111000000 : reciprocal = 1111111111111111;
        16'b1111101110111111 : reciprocal = 1111111111111111;
        16'b1111101110111110 : reciprocal = 1111111111111111;
        16'b1111101110111101 : reciprocal = 1111111111111111;
        16'b1111101110111100 : reciprocal = 1111111111111111;
        16'b1111101110111011 : reciprocal = 1111111111111111;
        16'b1111101110111010 : reciprocal = 1111111111111111;
        16'b1111101110111001 : reciprocal = 1111111111111111;
        16'b1111101110111000 : reciprocal = 1111111111111111;
        16'b1111101110110111 : reciprocal = 1111111111111111;
        16'b1111101110110110 : reciprocal = 1111111111111111;
        16'b1111101110110101 : reciprocal = 1111111111111111;
        16'b1111101110110100 : reciprocal = 1111111111111111;
        16'b1111101110110011 : reciprocal = 1111111111111111;
        16'b1111101110110010 : reciprocal = 1111111111111111;
        16'b1111101110110001 : reciprocal = 1111111111111111;
        16'b1111101110110000 : reciprocal = 1111111111111111;
        16'b1111101110101111 : reciprocal = 1111111111111111;
        16'b1111101110101110 : reciprocal = 1111111111111111;
        16'b1111101110101101 : reciprocal = 1111111111111111;
        16'b1111101110101100 : reciprocal = 1111111111111111;
        16'b1111101110101011 : reciprocal = 1111111111111111;
        16'b1111101110101010 : reciprocal = 1111111111111111;
        16'b1111101110101001 : reciprocal = 1111111111111111;
        16'b1111101110101000 : reciprocal = 1111111111111111;
        16'b1111101110100111 : reciprocal = 1111111111111111;
        16'b1111101110100110 : reciprocal = 1111111111111111;
        16'b1111101110100101 : reciprocal = 1111111111111111;
        16'b1111101110100100 : reciprocal = 1111111111111111;
        16'b1111101110100011 : reciprocal = 1111111111111111;
        16'b1111101110100010 : reciprocal = 1111111111111111;
        16'b1111101110100001 : reciprocal = 1111111111111111;
        16'b1111101110100000 : reciprocal = 1111111111111111;
        16'b1111101110011111 : reciprocal = 1111111111111111;
        16'b1111101110011110 : reciprocal = 1111111111111111;
        16'b1111101110011101 : reciprocal = 1111111111111111;
        16'b1111101110011100 : reciprocal = 1111111111111111;
        16'b1111101110011011 : reciprocal = 1111111111111111;
        16'b1111101110011010 : reciprocal = 1111111111111111;
        16'b1111101110011001 : reciprocal = 1111111111111111;
        16'b1111101110011000 : reciprocal = 1111111111111111;
        16'b1111101110010111 : reciprocal = 1111111111111111;
        16'b1111101110010110 : reciprocal = 1111111111111111;
        16'b1111101110010101 : reciprocal = 1111111111111111;
        16'b1111101110010100 : reciprocal = 1111111111111111;
        16'b1111101110010011 : reciprocal = 1111111111111111;
        16'b1111101110010010 : reciprocal = 1111111111111111;
        16'b1111101110010001 : reciprocal = 1111111111111111;
        16'b1111101110010000 : reciprocal = 1111111111111111;
        16'b1111101110001111 : reciprocal = 1111111111111111;
        16'b1111101110001110 : reciprocal = 1111111111111111;
        16'b1111101110001101 : reciprocal = 1111111111111111;
        16'b1111101110001100 : reciprocal = 1111111111111111;
        16'b1111101110001011 : reciprocal = 1111111111111111;
        16'b1111101110001010 : reciprocal = 1111111111111111;
        16'b1111101110001001 : reciprocal = 1111111111111111;
        16'b1111101110001000 : reciprocal = 1111111111111111;
        16'b1111101110000111 : reciprocal = 1111111111111111;
        16'b1111101110000110 : reciprocal = 1111111111111111;
        16'b1111101110000101 : reciprocal = 1111111111111111;
        16'b1111101110000100 : reciprocal = 1111111111111111;
        16'b1111101110000011 : reciprocal = 1111111111111111;
        16'b1111101110000010 : reciprocal = 1111111111111111;
        16'b1111101110000001 : reciprocal = 1111111111111111;
        16'b1111101110000000 : reciprocal = 1111111111111111;
        16'b1111101101111111 : reciprocal = 1111111111111111;
        16'b1111101101111110 : reciprocal = 1111111111111111;
        16'b1111101101111101 : reciprocal = 1111111111111111;
        16'b1111101101111100 : reciprocal = 1111111111111111;
        16'b1111101101111011 : reciprocal = 1111111111111111;
        16'b1111101101111010 : reciprocal = 1111111111111111;
        16'b1111101101111001 : reciprocal = 1111111111111111;
        16'b1111101101111000 : reciprocal = 1111111111111111;
        16'b1111101101110111 : reciprocal = 1111111111111111;
        16'b1111101101110110 : reciprocal = 1111111111111111;
        16'b1111101101110101 : reciprocal = 1111111111111111;
        16'b1111101101110100 : reciprocal = 1111111111111111;
        16'b1111101101110011 : reciprocal = 1111111111111111;
        16'b1111101101110010 : reciprocal = 1111111111111111;
        16'b1111101101110001 : reciprocal = 1111111111111111;
        16'b1111101101110000 : reciprocal = 1111111111111111;
        16'b1111101101101111 : reciprocal = 1111111111111111;
        16'b1111101101101110 : reciprocal = 1111111111111111;
        16'b1111101101101101 : reciprocal = 1111111111111111;
        16'b1111101101101100 : reciprocal = 1111111111111111;
        16'b1111101101101011 : reciprocal = 1111111111111111;
        16'b1111101101101010 : reciprocal = 1111111111111111;
        16'b1111101101101001 : reciprocal = 1111111111111111;
        16'b1111101101101000 : reciprocal = 1111111111111111;
        16'b1111101101100111 : reciprocal = 1111111111111111;
        16'b1111101101100110 : reciprocal = 1111111111111111;
        16'b1111101101100101 : reciprocal = 1111111111111111;
        16'b1111101101100100 : reciprocal = 1111111111111111;
        16'b1111101101100011 : reciprocal = 1111111111111111;
        16'b1111101101100010 : reciprocal = 1111111111111111;
        16'b1111101101100001 : reciprocal = 1111111111111111;
        16'b1111101101100000 : reciprocal = 1111111111111111;
        16'b1111101101011111 : reciprocal = 1111111111111111;
        16'b1111101101011110 : reciprocal = 1111111111111111;
        16'b1111101101011101 : reciprocal = 1111111111111111;
        16'b1111101101011100 : reciprocal = 1111111111111111;
        16'b1111101101011011 : reciprocal = 1111111111111111;
        16'b1111101101011010 : reciprocal = 1111111111111111;
        16'b1111101101011001 : reciprocal = 1111111111111111;
        16'b1111101101011000 : reciprocal = 1111111111111111;
        16'b1111101101010111 : reciprocal = 1111111111111111;
        16'b1111101101010110 : reciprocal = 1111111111111111;
        16'b1111101101010101 : reciprocal = 1111111111111111;
        16'b1111101101010100 : reciprocal = 1111111111111111;
        16'b1111101101010011 : reciprocal = 1111111111111111;
        16'b1111101101010010 : reciprocal = 1111111111111111;
        16'b1111101101010001 : reciprocal = 1111111111111111;
        16'b1111101101010000 : reciprocal = 1111111111111111;
        16'b1111101101001111 : reciprocal = 1111111111111111;
        16'b1111101101001110 : reciprocal = 1111111111111111;
        16'b1111101101001101 : reciprocal = 1111111111111111;
        16'b1111101101001100 : reciprocal = 1111111111111111;
        16'b1111101101001011 : reciprocal = 1111111111111111;
        16'b1111101101001010 : reciprocal = 1111111111111111;
        16'b1111101101001001 : reciprocal = 1111111111111111;
        16'b1111101101001000 : reciprocal = 1111111111111111;
        16'b1111101101000111 : reciprocal = 1111111111111111;
        16'b1111101101000110 : reciprocal = 1111111111111111;
        16'b1111101101000101 : reciprocal = 1111111111111111;
        16'b1111101101000100 : reciprocal = 1111111111111111;
        16'b1111101101000011 : reciprocal = 1111111111111111;
        16'b1111101101000010 : reciprocal = 1111111111111111;
        16'b1111101101000001 : reciprocal = 1111111111111111;
        16'b1111101101000000 : reciprocal = 1111111111111111;
        16'b1111101100111111 : reciprocal = 1111111111111111;
        16'b1111101100111110 : reciprocal = 1111111111111111;
        16'b1111101100111101 : reciprocal = 1111111111111111;
        16'b1111101100111100 : reciprocal = 1111111111111111;
        16'b1111101100111011 : reciprocal = 1111111111111111;
        16'b1111101100111010 : reciprocal = 1111111111111111;
        16'b1111101100111001 : reciprocal = 1111111111111111;
        16'b1111101100111000 : reciprocal = 1111111111111111;
        16'b1111101100110111 : reciprocal = 1111111111111111;
        16'b1111101100110110 : reciprocal = 1111111111111111;
        16'b1111101100110101 : reciprocal = 1111111111111111;
        16'b1111101100110100 : reciprocal = 1111111111111111;
        16'b1111101100110011 : reciprocal = 1111111111111111;
        16'b1111101100110010 : reciprocal = 1111111111111111;
        16'b1111101100110001 : reciprocal = 1111111111111111;
        16'b1111101100110000 : reciprocal = 1111111111111111;
        16'b1111101100101111 : reciprocal = 1111111111111111;
        16'b1111101100101110 : reciprocal = 1111111111111111;
        16'b1111101100101101 : reciprocal = 1111111111111111;
        16'b1111101100101100 : reciprocal = 1111111111111111;
        16'b1111101100101011 : reciprocal = 1111111111111111;
        16'b1111101100101010 : reciprocal = 1111111111111111;
        16'b1111101100101001 : reciprocal = 1111111111111111;
        16'b1111101100101000 : reciprocal = 1111111111111111;
        16'b1111101100100111 : reciprocal = 1111111111111111;
        16'b1111101100100110 : reciprocal = 1111111111111111;
        16'b1111101100100101 : reciprocal = 1111111111111111;
        16'b1111101100100100 : reciprocal = 1111111111111111;
        16'b1111101100100011 : reciprocal = 1111111111111111;
        16'b1111101100100010 : reciprocal = 1111111111111111;
        16'b1111101100100001 : reciprocal = 1111111111111111;
        16'b1111101100100000 : reciprocal = 1111111111111111;
        16'b1111101100011111 : reciprocal = 1111111111111111;
        16'b1111101100011110 : reciprocal = 1111111111111111;
        16'b1111101100011101 : reciprocal = 1111111111111111;
        16'b1111101100011100 : reciprocal = 1111111111111111;
        16'b1111101100011011 : reciprocal = 1111111111111111;
        16'b1111101100011010 : reciprocal = 1111111111111111;
        16'b1111101100011001 : reciprocal = 1111111111111111;
        16'b1111101100011000 : reciprocal = 1111111111111111;
        16'b1111101100010111 : reciprocal = 1111111111111111;
        16'b1111101100010110 : reciprocal = 1111111111111111;
        16'b1111101100010101 : reciprocal = 1111111111111111;
        16'b1111101100010100 : reciprocal = 1111111111111111;
        16'b1111101100010011 : reciprocal = 1111111111111111;
        16'b1111101100010010 : reciprocal = 1111111111111111;
        16'b1111101100010001 : reciprocal = 1111111111111111;
        16'b1111101100010000 : reciprocal = 1111111111111111;
        16'b1111101100001111 : reciprocal = 1111111111111111;
        16'b1111101100001110 : reciprocal = 1111111111111111;
        16'b1111101100001101 : reciprocal = 1111111111111111;
        16'b1111101100001100 : reciprocal = 1111111111111111;
        16'b1111101100001011 : reciprocal = 1111111111111111;
        16'b1111101100001010 : reciprocal = 1111111111111111;
        16'b1111101100001001 : reciprocal = 1111111111111111;
        16'b1111101100001000 : reciprocal = 1111111111111111;
        16'b1111101100000111 : reciprocal = 1111111111111111;
        16'b1111101100000110 : reciprocal = 1111111111111111;
        16'b1111101100000101 : reciprocal = 1111111111111111;
        16'b1111101100000100 : reciprocal = 1111111111111111;
        16'b1111101100000011 : reciprocal = 1111111111111111;
        16'b1111101100000010 : reciprocal = 1111111111111111;
        16'b1111101100000001 : reciprocal = 1111111111111111;
        16'b1111101100000000 : reciprocal = 1111111111111111;
        16'b1111101011111111 : reciprocal = 1111111111111111;
        16'b1111101011111110 : reciprocal = 1111111111111111;
        16'b1111101011111101 : reciprocal = 1111111111111111;
        16'b1111101011111100 : reciprocal = 1111111111111111;
        16'b1111101011111011 : reciprocal = 1111111111111111;
        16'b1111101011111010 : reciprocal = 1111111111111111;
        16'b1111101011111001 : reciprocal = 1111111111111111;
        16'b1111101011111000 : reciprocal = 1111111111111111;
        16'b1111101011110111 : reciprocal = 1111111111111111;
        16'b1111101011110110 : reciprocal = 1111111111111111;
        16'b1111101011110101 : reciprocal = 1111111111111111;
        16'b1111101011110100 : reciprocal = 1111111111111111;
        16'b1111101011110011 : reciprocal = 1111111111111111;
        16'b1111101011110010 : reciprocal = 1111111111111111;
        16'b1111101011110001 : reciprocal = 1111111111111111;
        16'b1111101011110000 : reciprocal = 1111111111111111;
        16'b1111101011101111 : reciprocal = 1111111111111111;
        16'b1111101011101110 : reciprocal = 1111111111111111;
        16'b1111101011101101 : reciprocal = 1111111111111111;
        16'b1111101011101100 : reciprocal = 1111111111111111;
        16'b1111101011101011 : reciprocal = 1111111111111111;
        16'b1111101011101010 : reciprocal = 1111111111111111;
        16'b1111101011101001 : reciprocal = 1111111111111111;
        16'b1111101011101000 : reciprocal = 1111111111111111;
        16'b1111101011100111 : reciprocal = 1111111111111111;
        16'b1111101011100110 : reciprocal = 1111111111111111;
        16'b1111101011100101 : reciprocal = 1111111111111111;
        16'b1111101011100100 : reciprocal = 1111111111111111;
        16'b1111101011100011 : reciprocal = 1111111111111111;
        16'b1111101011100010 : reciprocal = 1111111111111111;
        16'b1111101011100001 : reciprocal = 1111111111111111;
        16'b1111101011100000 : reciprocal = 1111111111111111;
        16'b1111101011011111 : reciprocal = 1111111111111111;
        16'b1111101011011110 : reciprocal = 1111111111111111;
        16'b1111101011011101 : reciprocal = 1111111111111111;
        16'b1111101011011100 : reciprocal = 1111111111111111;
        16'b1111101011011011 : reciprocal = 1111111111111111;
        16'b1111101011011010 : reciprocal = 1111111111111111;
        16'b1111101011011001 : reciprocal = 1111111111111111;
        16'b1111101011011000 : reciprocal = 1111111111111111;
        16'b1111101011010111 : reciprocal = 1111111111111111;
        16'b1111101011010110 : reciprocal = 1111111111111111;
        16'b1111101011010101 : reciprocal = 1111111111111111;
        16'b1111101011010100 : reciprocal = 1111111111111111;
        16'b1111101011010011 : reciprocal = 1111111111111111;
        16'b1111101011010010 : reciprocal = 1111111111111111;
        16'b1111101011010001 : reciprocal = 1111111111111111;
        16'b1111101011010000 : reciprocal = 1111111111111111;
        16'b1111101011001111 : reciprocal = 1111111111111111;
        16'b1111101011001110 : reciprocal = 1111111111111111;
        16'b1111101011001101 : reciprocal = 1111111111111111;
        16'b1111101011001100 : reciprocal = 1111111111111111;
        16'b1111101011001011 : reciprocal = 1111111111111111;
        16'b1111101011001010 : reciprocal = 1111111111111111;
        16'b1111101011001001 : reciprocal = 1111111111111111;
        16'b1111101011001000 : reciprocal = 1111111111111111;
        16'b1111101011000111 : reciprocal = 1111111111111111;
        16'b1111101011000110 : reciprocal = 1111111111111111;
        16'b1111101011000101 : reciprocal = 1111111111111111;
        16'b1111101011000100 : reciprocal = 1111111111111111;
        16'b1111101011000011 : reciprocal = 1111111111111111;
        16'b1111101011000010 : reciprocal = 1111111111111111;
        16'b1111101011000001 : reciprocal = 1111111111111111;
        16'b1111101011000000 : reciprocal = 1111111111111111;
        16'b1111101010111111 : reciprocal = 1111111111111111;
        16'b1111101010111110 : reciprocal = 1111111111111111;
        16'b1111101010111101 : reciprocal = 1111111111111111;
        16'b1111101010111100 : reciprocal = 1111111111111111;
        16'b1111101010111011 : reciprocal = 1111111111111111;
        16'b1111101010111010 : reciprocal = 1111111111111111;
        16'b1111101010111001 : reciprocal = 1111111111111111;
        16'b1111101010111000 : reciprocal = 1111111111111111;
        16'b1111101010110111 : reciprocal = 1111111111111111;
        16'b1111101010110110 : reciprocal = 1111111111111111;
        16'b1111101010110101 : reciprocal = 1111111111111111;
        16'b1111101010110100 : reciprocal = 1111111111111111;
        16'b1111101010110011 : reciprocal = 1111111111111111;
        16'b1111101010110010 : reciprocal = 1111111111111111;
        16'b1111101010110001 : reciprocal = 1111111111111111;
        16'b1111101010110000 : reciprocal = 1111111111111111;
        16'b1111101010101111 : reciprocal = 1111111111111111;
        16'b1111101010101110 : reciprocal = 1111111111111111;
        16'b1111101010101101 : reciprocal = 1111111111111111;
        16'b1111101010101100 : reciprocal = 1111111111111111;
        16'b1111101010101011 : reciprocal = 1111111111111111;
        16'b1111101010101010 : reciprocal = 1111111111111111;
        16'b1111101010101001 : reciprocal = 1111111111111111;
        16'b1111101010101000 : reciprocal = 1111111111111111;
        16'b1111101010100111 : reciprocal = 1111111111111111;
        16'b1111101010100110 : reciprocal = 1111111111111111;
        16'b1111101010100101 : reciprocal = 1111111111111111;
        16'b1111101010100100 : reciprocal = 1111111111111111;
        16'b1111101010100011 : reciprocal = 1111111111111111;
        16'b1111101010100010 : reciprocal = 1111111111111111;
        16'b1111101010100001 : reciprocal = 1111111111111111;
        16'b1111101010100000 : reciprocal = 1111111111111111;
        16'b1111101010011111 : reciprocal = 1111111111111111;
        16'b1111101010011110 : reciprocal = 1111111111111111;
        16'b1111101010011101 : reciprocal = 1111111111111111;
        16'b1111101010011100 : reciprocal = 1111111111111111;
        16'b1111101010011011 : reciprocal = 1111111111111111;
        16'b1111101010011010 : reciprocal = 1111111111111111;
        16'b1111101010011001 : reciprocal = 1111111111111111;
        16'b1111101010011000 : reciprocal = 1111111111111111;
        16'b1111101010010111 : reciprocal = 1111111111111111;
        16'b1111101010010110 : reciprocal = 1111111111111111;
        16'b1111101010010101 : reciprocal = 1111111111111111;
        16'b1111101010010100 : reciprocal = 1111111111111111;
        16'b1111101010010011 : reciprocal = 1111111111111111;
        16'b1111101010010010 : reciprocal = 1111111111111111;
        16'b1111101010010001 : reciprocal = 1111111111111111;
        16'b1111101010010000 : reciprocal = 1111111111111111;
        16'b1111101010001111 : reciprocal = 1111111111111111;
        16'b1111101010001110 : reciprocal = 1111111111111111;
        16'b1111101010001101 : reciprocal = 1111111111111111;
        16'b1111101010001100 : reciprocal = 1111111111111111;
        16'b1111101010001011 : reciprocal = 1111111111111111;
        16'b1111101010001010 : reciprocal = 1111111111111111;
        16'b1111101010001001 : reciprocal = 1111111111111111;
        16'b1111101010001000 : reciprocal = 1111111111111111;
        16'b1111101010000111 : reciprocal = 1111111111111111;
        16'b1111101010000110 : reciprocal = 1111111111111111;
        16'b1111101010000101 : reciprocal = 1111111111111111;
        16'b1111101010000100 : reciprocal = 1111111111111111;
        16'b1111101010000011 : reciprocal = 1111111111111111;
        16'b1111101010000010 : reciprocal = 1111111111111111;
        16'b1111101010000001 : reciprocal = 1111111111111111;
        16'b1111101010000000 : reciprocal = 1111111111111111;
        16'b1111101001111111 : reciprocal = 1111111111111111;
        16'b1111101001111110 : reciprocal = 1111111111111111;
        16'b1111101001111101 : reciprocal = 1111111111111111;
        16'b1111101001111100 : reciprocal = 1111111111111111;
        16'b1111101001111011 : reciprocal = 1111111111111111;
        16'b1111101001111010 : reciprocal = 1111111111111111;
        16'b1111101001111001 : reciprocal = 1111111111111111;
        16'b1111101001111000 : reciprocal = 1111111111111111;
        16'b1111101001110111 : reciprocal = 1111111111111111;
        16'b1111101001110110 : reciprocal = 1111111111111111;
        16'b1111101001110101 : reciprocal = 1111111111111111;
        16'b1111101001110100 : reciprocal = 1111111111111111;
        16'b1111101001110011 : reciprocal = 1111111111111111;
        16'b1111101001110010 : reciprocal = 1111111111111111;
        16'b1111101001110001 : reciprocal = 1111111111111111;
        16'b1111101001110000 : reciprocal = 1111111111111111;
        16'b1111101001101111 : reciprocal = 1111111111111111;
        16'b1111101001101110 : reciprocal = 1111111111111111;
        16'b1111101001101101 : reciprocal = 1111111111111111;
        16'b1111101001101100 : reciprocal = 1111111111111111;
        16'b1111101001101011 : reciprocal = 1111111111111111;
        16'b1111101001101010 : reciprocal = 1111111111111111;
        16'b1111101001101001 : reciprocal = 1111111111111111;
        16'b1111101001101000 : reciprocal = 1111111111111111;
        16'b1111101001100111 : reciprocal = 1111111111111111;
        16'b1111101001100110 : reciprocal = 1111111111111111;
        16'b1111101001100101 : reciprocal = 1111111111111111;
        16'b1111101001100100 : reciprocal = 1111111111111111;
        16'b1111101001100011 : reciprocal = 1111111111111111;
        16'b1111101001100010 : reciprocal = 1111111111111111;
        16'b1111101001100001 : reciprocal = 1111111111111111;
        16'b1111101001100000 : reciprocal = 1111111111111111;
        16'b1111101001011111 : reciprocal = 1111111111111111;
        16'b1111101001011110 : reciprocal = 1111111111111111;
        16'b1111101001011101 : reciprocal = 1111111111111111;
        16'b1111101001011100 : reciprocal = 1111111111111111;
        16'b1111101001011011 : reciprocal = 1111111111111111;
        16'b1111101001011010 : reciprocal = 1111111111111111;
        16'b1111101001011001 : reciprocal = 1111111111111111;
        16'b1111101001011000 : reciprocal = 1111111111111111;
        16'b1111101001010111 : reciprocal = 1111111111111111;
        16'b1111101001010110 : reciprocal = 1111111111111111;
        16'b1111101001010101 : reciprocal = 1111111111111111;
        16'b1111101001010100 : reciprocal = 1111111111111111;
        16'b1111101001010011 : reciprocal = 1111111111111111;
        16'b1111101001010010 : reciprocal = 1111111111111111;
        16'b1111101001010001 : reciprocal = 1111111111111111;
        16'b1111101001010000 : reciprocal = 1111111111111111;
        16'b1111101001001111 : reciprocal = 1111111111111111;
        16'b1111101001001110 : reciprocal = 1111111111111111;
        16'b1111101001001101 : reciprocal = 1111111111111111;
        16'b1111101001001100 : reciprocal = 1111111111111111;
        16'b1111101001001011 : reciprocal = 1111111111111111;
        16'b1111101001001010 : reciprocal = 1111111111111111;
        16'b1111101001001001 : reciprocal = 1111111111111111;
        16'b1111101001001000 : reciprocal = 1111111111111111;
        16'b1111101001000111 : reciprocal = 1111111111111111;
        16'b1111101001000110 : reciprocal = 1111111111111111;
        16'b1111101001000101 : reciprocal = 1111111111111111;
        16'b1111101001000100 : reciprocal = 1111111111111111;
        16'b1111101001000011 : reciprocal = 1111111111111111;
        16'b1111101001000010 : reciprocal = 1111111111111111;
        16'b1111101001000001 : reciprocal = 1111111111111111;
        16'b1111101001000000 : reciprocal = 1111111111111111;
        16'b1111101000111111 : reciprocal = 1111111111111111;
        16'b1111101000111110 : reciprocal = 1111111111111111;
        16'b1111101000111101 : reciprocal = 1111111111111111;
        16'b1111101000111100 : reciprocal = 1111111111111111;
        16'b1111101000111011 : reciprocal = 1111111111111111;
        16'b1111101000111010 : reciprocal = 1111111111111111;
        16'b1111101000111001 : reciprocal = 1111111111111111;
        16'b1111101000111000 : reciprocal = 1111111111111111;
        16'b1111101000110111 : reciprocal = 1111111111111111;
        16'b1111101000110110 : reciprocal = 1111111111111111;
        16'b1111101000110101 : reciprocal = 1111111111111111;
        16'b1111101000110100 : reciprocal = 1111111111111111;
        16'b1111101000110011 : reciprocal = 1111111111111111;
        16'b1111101000110010 : reciprocal = 1111111111111111;
        16'b1111101000110001 : reciprocal = 1111111111111111;
        16'b1111101000110000 : reciprocal = 1111111111111111;
        16'b1111101000101111 : reciprocal = 1111111111111111;
        16'b1111101000101110 : reciprocal = 1111111111111111;
        16'b1111101000101101 : reciprocal = 1111111111111111;
        16'b1111101000101100 : reciprocal = 1111111111111111;
        16'b1111101000101011 : reciprocal = 1111111111111111;
        16'b1111101000101010 : reciprocal = 1111111111111111;
        16'b1111101000101001 : reciprocal = 1111111111111111;
        16'b1111101000101000 : reciprocal = 1111111111111111;
        16'b1111101000100111 : reciprocal = 1111111111111111;
        16'b1111101000100110 : reciprocal = 1111111111111111;
        16'b1111101000100101 : reciprocal = 1111111111111111;
        16'b1111101000100100 : reciprocal = 1111111111111111;
        16'b1111101000100011 : reciprocal = 1111111111111111;
        16'b1111101000100010 : reciprocal = 1111111111111111;
        16'b1111101000100001 : reciprocal = 1111111111111111;
        16'b1111101000100000 : reciprocal = 1111111111111111;
        16'b1111101000011111 : reciprocal = 1111111111111111;
        16'b1111101000011110 : reciprocal = 1111111111111111;
        16'b1111101000011101 : reciprocal = 1111111111111111;
        16'b1111101000011100 : reciprocal = 1111111111111111;
        16'b1111101000011011 : reciprocal = 1111111111111111;
        16'b1111101000011010 : reciprocal = 1111111111111111;
        16'b1111101000011001 : reciprocal = 1111111111111111;
        16'b1111101000011000 : reciprocal = 1111111111111111;
        16'b1111101000010111 : reciprocal = 1111111111111111;
        16'b1111101000010110 : reciprocal = 1111111111111111;
        16'b1111101000010101 : reciprocal = 1111111111111111;
        16'b1111101000010100 : reciprocal = 1111111111111111;
        16'b1111101000010011 : reciprocal = 1111111111111111;
        16'b1111101000010010 : reciprocal = 1111111111111111;
        16'b1111101000010001 : reciprocal = 1111111111111111;
        16'b1111101000010000 : reciprocal = 1111111111111111;
        16'b1111101000001111 : reciprocal = 1111111111111111;
        16'b1111101000001110 : reciprocal = 1111111111111111;
        16'b1111101000001101 : reciprocal = 1111111111111111;
        16'b1111101000001100 : reciprocal = 1111111111111111;
        16'b1111101000001011 : reciprocal = 1111111111111111;
        16'b1111101000001010 : reciprocal = 1111111111111111;
        16'b1111101000001001 : reciprocal = 1111111111111111;
        16'b1111101000001000 : reciprocal = 1111111111111111;
        16'b1111101000000111 : reciprocal = 1111111111111111;
        16'b1111101000000110 : reciprocal = 1111111111111111;
        16'b1111101000000101 : reciprocal = 1111111111111111;
        16'b1111101000000100 : reciprocal = 1111111111111111;
        16'b1111101000000011 : reciprocal = 1111111111111111;
        16'b1111101000000010 : reciprocal = 1111111111111111;
        16'b1111101000000001 : reciprocal = 1111111111111111;
        16'b1111101000000000 : reciprocal = 1111111111111111;
        16'b1111100111111111 : reciprocal = 1111111111111111;
        16'b1111100111111110 : reciprocal = 1111111111111111;
        16'b1111100111111101 : reciprocal = 1111111111111111;
        16'b1111100111111100 : reciprocal = 1111111111111111;
        16'b1111100111111011 : reciprocal = 1111111111111111;
        16'b1111100111111010 : reciprocal = 1111111111111111;
        16'b1111100111111001 : reciprocal = 1111111111111111;
        16'b1111100111111000 : reciprocal = 1111111111111111;
        16'b1111100111110111 : reciprocal = 1111111111111111;
        16'b1111100111110110 : reciprocal = 1111111111111111;
        16'b1111100111110101 : reciprocal = 1111111111111111;
        16'b1111100111110100 : reciprocal = 1111111111111111;
        16'b1111100111110011 : reciprocal = 1111111111111111;
        16'b1111100111110010 : reciprocal = 1111111111111111;
        16'b1111100111110001 : reciprocal = 1111111111111111;
        16'b1111100111110000 : reciprocal = 1111111111111111;
        16'b1111100111101111 : reciprocal = 1111111111111111;
        16'b1111100111101110 : reciprocal = 1111111111111111;
        16'b1111100111101101 : reciprocal = 1111111111111111;
        16'b1111100111101100 : reciprocal = 1111111111111111;
        16'b1111100111101011 : reciprocal = 1111111111111111;
        16'b1111100111101010 : reciprocal = 1111111111111111;
        16'b1111100111101001 : reciprocal = 1111111111111111;
        16'b1111100111101000 : reciprocal = 1111111111111111;
        16'b1111100111100111 : reciprocal = 1111111111111111;
        16'b1111100111100110 : reciprocal = 1111111111111111;
        16'b1111100111100101 : reciprocal = 1111111111111111;
        16'b1111100111100100 : reciprocal = 1111111111111111;
        16'b1111100111100011 : reciprocal = 1111111111111111;
        16'b1111100111100010 : reciprocal = 1111111111111111;
        16'b1111100111100001 : reciprocal = 1111111111111111;
        16'b1111100111100000 : reciprocal = 1111111111111111;
        16'b1111100111011111 : reciprocal = 1111111111111111;
        16'b1111100111011110 : reciprocal = 1111111111111111;
        16'b1111100111011101 : reciprocal = 1111111111111111;
        16'b1111100111011100 : reciprocal = 1111111111111111;
        16'b1111100111011011 : reciprocal = 1111111111111111;
        16'b1111100111011010 : reciprocal = 1111111111111111;
        16'b1111100111011001 : reciprocal = 1111111111111111;
        16'b1111100111011000 : reciprocal = 1111111111111111;
        16'b1111100111010111 : reciprocal = 1111111111111111;
        16'b1111100111010110 : reciprocal = 1111111111111111;
        16'b1111100111010101 : reciprocal = 1111111111111111;
        16'b1111100111010100 : reciprocal = 1111111111111111;
        16'b1111100111010011 : reciprocal = 1111111111111111;
        16'b1111100111010010 : reciprocal = 1111111111111111;
        16'b1111100111010001 : reciprocal = 1111111111111111;
        16'b1111100111010000 : reciprocal = 1111111111111111;
        16'b1111100111001111 : reciprocal = 1111111111111111;
        16'b1111100111001110 : reciprocal = 1111111111111111;
        16'b1111100111001101 : reciprocal = 1111111111111111;
        16'b1111100111001100 : reciprocal = 1111111111111111;
        16'b1111100111001011 : reciprocal = 1111111111111111;
        16'b1111100111001010 : reciprocal = 1111111111111111;
        16'b1111100111001001 : reciprocal = 1111111111111111;
        16'b1111100111001000 : reciprocal = 1111111111111111;
        16'b1111100111000111 : reciprocal = 1111111111111111;
        16'b1111100111000110 : reciprocal = 1111111111111111;
        16'b1111100111000101 : reciprocal = 1111111111111111;
        16'b1111100111000100 : reciprocal = 1111111111111111;
        16'b1111100111000011 : reciprocal = 1111111111111111;
        16'b1111100111000010 : reciprocal = 1111111111111111;
        16'b1111100111000001 : reciprocal = 1111111111111111;
        16'b1111100111000000 : reciprocal = 1111111111111111;
        16'b1111100110111111 : reciprocal = 1111111111111111;
        16'b1111100110111110 : reciprocal = 1111111111111111;
        16'b1111100110111101 : reciprocal = 1111111111111111;
        16'b1111100110111100 : reciprocal = 1111111111111111;
        16'b1111100110111011 : reciprocal = 1111111111111111;
        16'b1111100110111010 : reciprocal = 1111111111111111;
        16'b1111100110111001 : reciprocal = 1111111111111111;
        16'b1111100110111000 : reciprocal = 1111111111111111;
        16'b1111100110110111 : reciprocal = 1111111111111111;
        16'b1111100110110110 : reciprocal = 1111111111111111;
        16'b1111100110110101 : reciprocal = 1111111111111111;
        16'b1111100110110100 : reciprocal = 1111111111111111;
        16'b1111100110110011 : reciprocal = 1111111111111111;
        16'b1111100110110010 : reciprocal = 1111111111111111;
        16'b1111100110110001 : reciprocal = 1111111111111111;
        16'b1111100110110000 : reciprocal = 1111111111111111;
        16'b1111100110101111 : reciprocal = 1111111111111111;
        16'b1111100110101110 : reciprocal = 1111111111111111;
        16'b1111100110101101 : reciprocal = 1111111111111111;
        16'b1111100110101100 : reciprocal = 1111111111111111;
        16'b1111100110101011 : reciprocal = 1111111111111111;
        16'b1111100110101010 : reciprocal = 1111111111111111;
        16'b1111100110101001 : reciprocal = 1111111111111111;
        16'b1111100110101000 : reciprocal = 1111111111111111;
        16'b1111100110100111 : reciprocal = 1111111111111111;
        16'b1111100110100110 : reciprocal = 1111111111111111;
        16'b1111100110100101 : reciprocal = 1111111111111111;
        16'b1111100110100100 : reciprocal = 1111111111111111;
        16'b1111100110100011 : reciprocal = 1111111111111111;
        16'b1111100110100010 : reciprocal = 1111111111111111;
        16'b1111100110100001 : reciprocal = 1111111111111111;
        16'b1111100110100000 : reciprocal = 1111111111111111;
        16'b1111100110011111 : reciprocal = 1111111111111111;
        16'b1111100110011110 : reciprocal = 1111111111111111;
        16'b1111100110011101 : reciprocal = 1111111111111111;
        16'b1111100110011100 : reciprocal = 1111111111111111;
        16'b1111100110011011 : reciprocal = 1111111111111111;
        16'b1111100110011010 : reciprocal = 1111111111111111;
        16'b1111100110011001 : reciprocal = 1111111111111111;
        16'b1111100110011000 : reciprocal = 1111111111111111;
        16'b1111100110010111 : reciprocal = 1111111111111111;
        16'b1111100110010110 : reciprocal = 1111111111111111;
        16'b1111100110010101 : reciprocal = 1111111111111111;
        16'b1111100110010100 : reciprocal = 1111111111111111;
        16'b1111100110010011 : reciprocal = 1111111111111111;
        16'b1111100110010010 : reciprocal = 1111111111111111;
        16'b1111100110010001 : reciprocal = 1111111111111111;
        16'b1111100110010000 : reciprocal = 1111111111111111;
        16'b1111100110001111 : reciprocal = 1111111111111111;
        16'b1111100110001110 : reciprocal = 1111111111111111;
        16'b1111100110001101 : reciprocal = 1111111111111111;
        16'b1111100110001100 : reciprocal = 1111111111111111;
        16'b1111100110001011 : reciprocal = 1111111111111111;
        16'b1111100110001010 : reciprocal = 1111111111111111;
        16'b1111100110001001 : reciprocal = 1111111111111111;
        16'b1111100110001000 : reciprocal = 1111111111111111;
        16'b1111100110000111 : reciprocal = 1111111111111111;
        16'b1111100110000110 : reciprocal = 1111111111111111;
        16'b1111100110000101 : reciprocal = 1111111111111111;
        16'b1111100110000100 : reciprocal = 1111111111111111;
        16'b1111100110000011 : reciprocal = 1111111111111111;
        16'b1111100110000010 : reciprocal = 1111111111111111;
        16'b1111100110000001 : reciprocal = 1111111111111111;
        16'b1111100110000000 : reciprocal = 1111111111111111;
        16'b1111100101111111 : reciprocal = 1111111111111111;
        16'b1111100101111110 : reciprocal = 1111111111111111;
        16'b1111100101111101 : reciprocal = 1111111111111111;
        16'b1111100101111100 : reciprocal = 1111111111111111;
        16'b1111100101111011 : reciprocal = 1111111111111111;
        16'b1111100101111010 : reciprocal = 1111111111111111;
        16'b1111100101111001 : reciprocal = 1111111111111111;
        16'b1111100101111000 : reciprocal = 1111111111111111;
        16'b1111100101110111 : reciprocal = 1111111111111111;
        16'b1111100101110110 : reciprocal = 1111111111111111;
        16'b1111100101110101 : reciprocal = 1111111111111111;
        16'b1111100101110100 : reciprocal = 1111111111111111;
        16'b1111100101110011 : reciprocal = 1111111111111111;
        16'b1111100101110010 : reciprocal = 1111111111111111;
        16'b1111100101110001 : reciprocal = 1111111111111111;
        16'b1111100101110000 : reciprocal = 1111111111111111;
        16'b1111100101101111 : reciprocal = 1111111111111111;
        16'b1111100101101110 : reciprocal = 1111111111111111;
        16'b1111100101101101 : reciprocal = 1111111111111111;
        16'b1111100101101100 : reciprocal = 1111111111111111;
        16'b1111100101101011 : reciprocal = 1111111111111111;
        16'b1111100101101010 : reciprocal = 1111111111111111;
        16'b1111100101101001 : reciprocal = 1111111111111111;
        16'b1111100101101000 : reciprocal = 1111111111111111;
        16'b1111100101100111 : reciprocal = 1111111111111111;
        16'b1111100101100110 : reciprocal = 1111111111111111;
        16'b1111100101100101 : reciprocal = 1111111111111111;
        16'b1111100101100100 : reciprocal = 1111111111111111;
        16'b1111100101100011 : reciprocal = 1111111111111111;
        16'b1111100101100010 : reciprocal = 1111111111111111;
        16'b1111100101100001 : reciprocal = 1111111111111111;
        16'b1111100101100000 : reciprocal = 1111111111111111;
        16'b1111100101011111 : reciprocal = 1111111111111111;
        16'b1111100101011110 : reciprocal = 1111111111111111;
        16'b1111100101011101 : reciprocal = 1111111111111111;
        16'b1111100101011100 : reciprocal = 1111111111111111;
        16'b1111100101011011 : reciprocal = 1111111111111111;
        16'b1111100101011010 : reciprocal = 1111111111111111;
        16'b1111100101011001 : reciprocal = 1111111111111111;
        16'b1111100101011000 : reciprocal = 1111111111111111;
        16'b1111100101010111 : reciprocal = 1111111111111111;
        16'b1111100101010110 : reciprocal = 1111111111111111;
        16'b1111100101010101 : reciprocal = 1111111111111111;
        16'b1111100101010100 : reciprocal = 1111111111111111;
        16'b1111100101010011 : reciprocal = 1111111111111111;
        16'b1111100101010010 : reciprocal = 1111111111111111;
        16'b1111100101010001 : reciprocal = 1111111111111111;
        16'b1111100101010000 : reciprocal = 1111111111111111;
        16'b1111100101001111 : reciprocal = 1111111111111111;
        16'b1111100101001110 : reciprocal = 1111111111111111;
        16'b1111100101001101 : reciprocal = 1111111111111111;
        16'b1111100101001100 : reciprocal = 1111111111111111;
        16'b1111100101001011 : reciprocal = 1111111111111111;
        16'b1111100101001010 : reciprocal = 1111111111111111;
        16'b1111100101001001 : reciprocal = 1111111111111111;
        16'b1111100101001000 : reciprocal = 1111111111111111;
        16'b1111100101000111 : reciprocal = 1111111111111111;
        16'b1111100101000110 : reciprocal = 1111111111111111;
        16'b1111100101000101 : reciprocal = 1111111111111111;
        16'b1111100101000100 : reciprocal = 1111111111111111;
        16'b1111100101000011 : reciprocal = 1111111111111111;
        16'b1111100101000010 : reciprocal = 1111111111111111;
        16'b1111100101000001 : reciprocal = 1111111111111111;
        16'b1111100101000000 : reciprocal = 1111111111111111;
        16'b1111100100111111 : reciprocal = 1111111111111111;
        16'b1111100100111110 : reciprocal = 1111111111111111;
        16'b1111100100111101 : reciprocal = 1111111111111111;
        16'b1111100100111100 : reciprocal = 1111111111111111;
        16'b1111100100111011 : reciprocal = 1111111111111111;
        16'b1111100100111010 : reciprocal = 1111111111111111;
        16'b1111100100111001 : reciprocal = 1111111111111111;
        16'b1111100100111000 : reciprocal = 1111111111111111;
        16'b1111100100110111 : reciprocal = 1111111111111111;
        16'b1111100100110110 : reciprocal = 1111111111111111;
        16'b1111100100110101 : reciprocal = 1111111111111111;
        16'b1111100100110100 : reciprocal = 1111111111111111;
        16'b1111100100110011 : reciprocal = 1111111111111111;
        16'b1111100100110010 : reciprocal = 1111111111111111;
        16'b1111100100110001 : reciprocal = 1111111111111111;
        16'b1111100100110000 : reciprocal = 1111111111111111;
        16'b1111100100101111 : reciprocal = 1111111111111111;
        16'b1111100100101110 : reciprocal = 1111111111111111;
        16'b1111100100101101 : reciprocal = 1111111111111111;
        16'b1111100100101100 : reciprocal = 1111111111111111;
        16'b1111100100101011 : reciprocal = 1111111111111111;
        16'b1111100100101010 : reciprocal = 1111111111111111;
        16'b1111100100101001 : reciprocal = 1111111111111111;
        16'b1111100100101000 : reciprocal = 1111111111111111;
        16'b1111100100100111 : reciprocal = 1111111111111111;
        16'b1111100100100110 : reciprocal = 1111111111111111;
        16'b1111100100100101 : reciprocal = 1111111111111111;
        16'b1111100100100100 : reciprocal = 1111111111111111;
        16'b1111100100100011 : reciprocal = 1111111111111111;
        16'b1111100100100010 : reciprocal = 1111111111111111;
        16'b1111100100100001 : reciprocal = 1111111111111111;
        16'b1111100100100000 : reciprocal = 1111111111111111;
        16'b1111100100011111 : reciprocal = 1111111111111111;
        16'b1111100100011110 : reciprocal = 1111111111111111;
        16'b1111100100011101 : reciprocal = 1111111111111111;
        16'b1111100100011100 : reciprocal = 1111111111111111;
        16'b1111100100011011 : reciprocal = 1111111111111111;
        16'b1111100100011010 : reciprocal = 1111111111111111;
        16'b1111100100011001 : reciprocal = 1111111111111111;
        16'b1111100100011000 : reciprocal = 1111111111111111;
        16'b1111100100010111 : reciprocal = 1111111111111111;
        16'b1111100100010110 : reciprocal = 1111111111111111;
        16'b1111100100010101 : reciprocal = 1111111111111111;
        16'b1111100100010100 : reciprocal = 1111111111111111;
        16'b1111100100010011 : reciprocal = 1111111111111111;
        16'b1111100100010010 : reciprocal = 1111111111111111;
        16'b1111100100010001 : reciprocal = 1111111111111111;
        16'b1111100100010000 : reciprocal = 1111111111111111;
        16'b1111100100001111 : reciprocal = 1111111111111111;
        16'b1111100100001110 : reciprocal = 1111111111111111;
        16'b1111100100001101 : reciprocal = 1111111111111111;
        16'b1111100100001100 : reciprocal = 1111111111111111;
        16'b1111100100001011 : reciprocal = 1111111111111111;
        16'b1111100100001010 : reciprocal = 1111111111111111;
        16'b1111100100001001 : reciprocal = 1111111111111111;
        16'b1111100100001000 : reciprocal = 1111111111111111;
        16'b1111100100000111 : reciprocal = 1111111111111111;
        16'b1111100100000110 : reciprocal = 1111111111111111;
        16'b1111100100000101 : reciprocal = 1111111111111111;
        16'b1111100100000100 : reciprocal = 1111111111111111;
        16'b1111100100000011 : reciprocal = 1111111111111111;
        16'b1111100100000010 : reciprocal = 1111111111111111;
        16'b1111100100000001 : reciprocal = 1111111111111111;
        16'b1111100100000000 : reciprocal = 1111111111111111;
        16'b1111100011111111 : reciprocal = 1111111111111111;
        16'b1111100011111110 : reciprocal = 1111111111111111;
        16'b1111100011111101 : reciprocal = 1111111111111111;
        16'b1111100011111100 : reciprocal = 1111111111111111;
        16'b1111100011111011 : reciprocal = 1111111111111111;
        16'b1111100011111010 : reciprocal = 1111111111111111;
        16'b1111100011111001 : reciprocal = 1111111111111111;
        16'b1111100011111000 : reciprocal = 1111111111111111;
        16'b1111100011110111 : reciprocal = 1111111111111111;
        16'b1111100011110110 : reciprocal = 1111111111111111;
        16'b1111100011110101 : reciprocal = 1111111111111111;
        16'b1111100011110100 : reciprocal = 1111111111111111;
        16'b1111100011110011 : reciprocal = 1111111111111111;
        16'b1111100011110010 : reciprocal = 1111111111111111;
        16'b1111100011110001 : reciprocal = 1111111111111111;
        16'b1111100011110000 : reciprocal = 1111111111111111;
        16'b1111100011101111 : reciprocal = 1111111111111111;
        16'b1111100011101110 : reciprocal = 1111111111111111;
        16'b1111100011101101 : reciprocal = 1111111111111111;
        16'b1111100011101100 : reciprocal = 1111111111111111;
        16'b1111100011101011 : reciprocal = 1111111111111111;
        16'b1111100011101010 : reciprocal = 1111111111111111;
        16'b1111100011101001 : reciprocal = 1111111111111111;
        16'b1111100011101000 : reciprocal = 1111111111111111;
        16'b1111100011100111 : reciprocal = 1111111111111111;
        16'b1111100011100110 : reciprocal = 1111111111111111;
        16'b1111100011100101 : reciprocal = 1111111111111111;
        16'b1111100011100100 : reciprocal = 1111111111111111;
        16'b1111100011100011 : reciprocal = 1111111111111111;
        16'b1111100011100010 : reciprocal = 1111111111111111;
        16'b1111100011100001 : reciprocal = 1111111111111111;
        16'b1111100011100000 : reciprocal = 1111111111111111;
        16'b1111100011011111 : reciprocal = 1111111111111111;
        16'b1111100011011110 : reciprocal = 1111111111111111;
        16'b1111100011011101 : reciprocal = 1111111111111111;
        16'b1111100011011100 : reciprocal = 1111111111111111;
        16'b1111100011011011 : reciprocal = 1111111111111111;
        16'b1111100011011010 : reciprocal = 1111111111111111;
        16'b1111100011011001 : reciprocal = 1111111111111111;
        16'b1111100011011000 : reciprocal = 1111111111111111;
        16'b1111100011010111 : reciprocal = 1111111111111111;
        16'b1111100011010110 : reciprocal = 1111111111111111;
        16'b1111100011010101 : reciprocal = 1111111111111111;
        16'b1111100011010100 : reciprocal = 1111111111111111;
        16'b1111100011010011 : reciprocal = 1111111111111111;
        16'b1111100011010010 : reciprocal = 1111111111111111;
        16'b1111100011010001 : reciprocal = 1111111111111111;
        16'b1111100011010000 : reciprocal = 1111111111111111;
        16'b1111100011001111 : reciprocal = 1111111111111111;
        16'b1111100011001110 : reciprocal = 1111111111111111;
        16'b1111100011001101 : reciprocal = 1111111111111111;
        16'b1111100011001100 : reciprocal = 1111111111111111;
        16'b1111100011001011 : reciprocal = 1111111111111111;
        16'b1111100011001010 : reciprocal = 1111111111111111;
        16'b1111100011001001 : reciprocal = 1111111111111111;
        16'b1111100011001000 : reciprocal = 1111111111111111;
        16'b1111100011000111 : reciprocal = 1111111111111111;
        16'b1111100011000110 : reciprocal = 1111111111111111;
        16'b1111100011000101 : reciprocal = 1111111111111111;
        16'b1111100011000100 : reciprocal = 1111111111111111;
        16'b1111100011000011 : reciprocal = 1111111111111111;
        16'b1111100011000010 : reciprocal = 1111111111111111;
        16'b1111100011000001 : reciprocal = 1111111111111111;
        16'b1111100011000000 : reciprocal = 1111111111111111;
        16'b1111100010111111 : reciprocal = 1111111111111111;
        16'b1111100010111110 : reciprocal = 1111111111111111;
        16'b1111100010111101 : reciprocal = 1111111111111111;
        16'b1111100010111100 : reciprocal = 1111111111111111;
        16'b1111100010111011 : reciprocal = 1111111111111111;
        16'b1111100010111010 : reciprocal = 1111111111111111;
        16'b1111100010111001 : reciprocal = 1111111111111111;
        16'b1111100010111000 : reciprocal = 1111111111111111;
        16'b1111100010110111 : reciprocal = 1111111111111111;
        16'b1111100010110110 : reciprocal = 1111111111111111;
        16'b1111100010110101 : reciprocal = 1111111111111111;
        16'b1111100010110100 : reciprocal = 1111111111111111;
        16'b1111100010110011 : reciprocal = 1111111111111111;
        16'b1111100010110010 : reciprocal = 1111111111111111;
        16'b1111100010110001 : reciprocal = 1111111111111111;
        16'b1111100010110000 : reciprocal = 1111111111111111;
        16'b1111100010101111 : reciprocal = 1111111111111111;
        16'b1111100010101110 : reciprocal = 1111111111111111;
        16'b1111100010101101 : reciprocal = 1111111111111111;
        16'b1111100010101100 : reciprocal = 1111111111111111;
        16'b1111100010101011 : reciprocal = 1111111111111111;
        16'b1111100010101010 : reciprocal = 1111111111111111;
        16'b1111100010101001 : reciprocal = 1111111111111111;
        16'b1111100010101000 : reciprocal = 1111111111111111;
        16'b1111100010100111 : reciprocal = 1111111111111111;
        16'b1111100010100110 : reciprocal = 1111111111111111;
        16'b1111100010100101 : reciprocal = 1111111111111111;
        16'b1111100010100100 : reciprocal = 1111111111111111;
        16'b1111100010100011 : reciprocal = 1111111111111111;
        16'b1111100010100010 : reciprocal = 1111111111111111;
        16'b1111100010100001 : reciprocal = 1111111111111111;
        16'b1111100010100000 : reciprocal = 1111111111111111;
        16'b1111100010011111 : reciprocal = 1111111111111111;
        16'b1111100010011110 : reciprocal = 1111111111111111;
        16'b1111100010011101 : reciprocal = 1111111111111111;
        16'b1111100010011100 : reciprocal = 1111111111111111;
        16'b1111100010011011 : reciprocal = 1111111111111111;
        16'b1111100010011010 : reciprocal = 1111111111111111;
        16'b1111100010011001 : reciprocal = 1111111111111111;
        16'b1111100010011000 : reciprocal = 1111111111111111;
        16'b1111100010010111 : reciprocal = 1111111111111111;
        16'b1111100010010110 : reciprocal = 1111111111111111;
        16'b1111100010010101 : reciprocal = 1111111111111111;
        16'b1111100010010100 : reciprocal = 1111111111111111;
        16'b1111100010010011 : reciprocal = 1111111111111111;
        16'b1111100010010010 : reciprocal = 1111111111111111;
        16'b1111100010010001 : reciprocal = 1111111111111111;
        16'b1111100010010000 : reciprocal = 1111111111111111;
        16'b1111100010001111 : reciprocal = 1111111111111111;
        16'b1111100010001110 : reciprocal = 1111111111111111;
        16'b1111100010001101 : reciprocal = 1111111111111111;
        16'b1111100010001100 : reciprocal = 1111111111111111;
        16'b1111100010001011 : reciprocal = 1111111111111111;
        16'b1111100010001010 : reciprocal = 1111111111111111;
        16'b1111100010001001 : reciprocal = 1111111111111111;
        16'b1111100010001000 : reciprocal = 1111111111111111;
        16'b1111100010000111 : reciprocal = 1111111111111111;
        16'b1111100010000110 : reciprocal = 1111111111111111;
        16'b1111100010000101 : reciprocal = 1111111111111111;
        16'b1111100010000100 : reciprocal = 1111111111111111;
        16'b1111100010000011 : reciprocal = 1111111111111111;
        16'b1111100010000010 : reciprocal = 1111111111111111;
        16'b1111100010000001 : reciprocal = 1111111111111111;
        16'b1111100010000000 : reciprocal = 1111111111111111;
        16'b1111100001111111 : reciprocal = 1111111111111111;
        16'b1111100001111110 : reciprocal = 1111111111111111;
        16'b1111100001111101 : reciprocal = 1111111111111111;
        16'b1111100001111100 : reciprocal = 1111111111111111;
        16'b1111100001111011 : reciprocal = 1111111111111111;
        16'b1111100001111010 : reciprocal = 1111111111111111;
        16'b1111100001111001 : reciprocal = 1111111111111111;
        16'b1111100001111000 : reciprocal = 1111111111111111;
        16'b1111100001110111 : reciprocal = 1111111111111111;
        16'b1111100001110110 : reciprocal = 1111111111111111;
        16'b1111100001110101 : reciprocal = 1111111111111111;
        16'b1111100001110100 : reciprocal = 1111111111111111;
        16'b1111100001110011 : reciprocal = 1111111111111111;
        16'b1111100001110010 : reciprocal = 1111111111111111;
        16'b1111100001110001 : reciprocal = 1111111111111111;
        16'b1111100001110000 : reciprocal = 1111111111111111;
        16'b1111100001101111 : reciprocal = 1111111111111111;
        16'b1111100001101110 : reciprocal = 1111111111111111;
        16'b1111100001101101 : reciprocal = 1111111111111111;
        16'b1111100001101100 : reciprocal = 1111111111111111;
        16'b1111100001101011 : reciprocal = 1111111111111111;
        16'b1111100001101010 : reciprocal = 1111111111111111;
        16'b1111100001101001 : reciprocal = 1111111111111111;
        16'b1111100001101000 : reciprocal = 1111111111111111;
        16'b1111100001100111 : reciprocal = 1111111111111111;
        16'b1111100001100110 : reciprocal = 1111111111111111;
        16'b1111100001100101 : reciprocal = 1111111111111111;
        16'b1111100001100100 : reciprocal = 1111111111111111;
        16'b1111100001100011 : reciprocal = 1111111111111111;
        16'b1111100001100010 : reciprocal = 1111111111111111;
        16'b1111100001100001 : reciprocal = 1111111111111111;
        16'b1111100001100000 : reciprocal = 1111111111111111;
        16'b1111100001011111 : reciprocal = 1111111111111111;
        16'b1111100001011110 : reciprocal = 1111111111111111;
        16'b1111100001011101 : reciprocal = 1111111111111111;
        16'b1111100001011100 : reciprocal = 1111111111111111;
        16'b1111100001011011 : reciprocal = 1111111111111111;
        16'b1111100001011010 : reciprocal = 1111111111111111;
        16'b1111100001011001 : reciprocal = 1111111111111111;
        16'b1111100001011000 : reciprocal = 1111111111111111;
        16'b1111100001010111 : reciprocal = 1111111111111111;
        16'b1111100001010110 : reciprocal = 1111111111111111;
        16'b1111100001010101 : reciprocal = 1111111111111111;
        16'b1111100001010100 : reciprocal = 1111111111111111;
        16'b1111100001010011 : reciprocal = 1111111111111111;
        16'b1111100001010010 : reciprocal = 1111111111111111;
        16'b1111100001010001 : reciprocal = 1111111111111111;
        16'b1111100001010000 : reciprocal = 1111111111111111;
        16'b1111100001001111 : reciprocal = 1111111111111111;
        16'b1111100001001110 : reciprocal = 1111111111111111;
        16'b1111100001001101 : reciprocal = 1111111111111111;
        16'b1111100001001100 : reciprocal = 1111111111111111;
        16'b1111100001001011 : reciprocal = 1111111111111111;
        16'b1111100001001010 : reciprocal = 1111111111111111;
        16'b1111100001001001 : reciprocal = 1111111111111111;
        16'b1111100001001000 : reciprocal = 1111111111111111;
        16'b1111100001000111 : reciprocal = 1111111111111111;
        16'b1111100001000110 : reciprocal = 1111111111111111;
        16'b1111100001000101 : reciprocal = 1111111111111111;
        16'b1111100001000100 : reciprocal = 1111111111111111;
        16'b1111100001000011 : reciprocal = 1111111111111111;
        16'b1111100001000010 : reciprocal = 1111111111111111;
        16'b1111100001000001 : reciprocal = 1111111111111111;
        16'b1111100001000000 : reciprocal = 1111111111111111;
        16'b1111100000111111 : reciprocal = 1111111111111111;
        16'b1111100000111110 : reciprocal = 1111111111111111;
        16'b1111100000111101 : reciprocal = 1111111111111111;
        16'b1111100000111100 : reciprocal = 1111111111111111;
        16'b1111100000111011 : reciprocal = 1111111111111111;
        16'b1111100000111010 : reciprocal = 1111111111111111;
        16'b1111100000111001 : reciprocal = 1111111111111111;
        16'b1111100000111000 : reciprocal = 1111111111111111;
        16'b1111100000110111 : reciprocal = 1111111111111111;
        16'b1111100000110110 : reciprocal = 1111111111111111;
        16'b1111100000110101 : reciprocal = 1111111111111111;
        16'b1111100000110100 : reciprocal = 1111111111111111;
        16'b1111100000110011 : reciprocal = 1111111111111111;
        16'b1111100000110010 : reciprocal = 1111111111111111;
        16'b1111100000110001 : reciprocal = 1111111111111111;
        16'b1111100000110000 : reciprocal = 1111111111111111;
        16'b1111100000101111 : reciprocal = 1111111111111111;
        16'b1111100000101110 : reciprocal = 1111111111111111;
        16'b1111100000101101 : reciprocal = 1111111111111111;
        16'b1111100000101100 : reciprocal = 1111111111111111;
        16'b1111100000101011 : reciprocal = 1111111111111111;
        16'b1111100000101010 : reciprocal = 1111111111111111;
        16'b1111100000101001 : reciprocal = 1111111111111111;
        16'b1111100000101000 : reciprocal = 1111111111111111;
        16'b1111100000100111 : reciprocal = 1111111111111111;
        16'b1111100000100110 : reciprocal = 1111111111111111;
        16'b1111100000100101 : reciprocal = 1111111111111111;
        16'b1111100000100100 : reciprocal = 1111111111111111;
        16'b1111100000100011 : reciprocal = 1111111111111111;
        16'b1111100000100010 : reciprocal = 1111111111111111;
        16'b1111100000100001 : reciprocal = 1111111111111111;
        16'b1111100000100000 : reciprocal = 1111111111111111;
        16'b1111100000011111 : reciprocal = 1111111111111111;
        16'b1111100000011110 : reciprocal = 1111111111111111;
        16'b1111100000011101 : reciprocal = 1111111111111111;
        16'b1111100000011100 : reciprocal = 1111111111111111;
        16'b1111100000011011 : reciprocal = 1111111111111111;
        16'b1111100000011010 : reciprocal = 1111111111111111;
        16'b1111100000011001 : reciprocal = 1111111111111111;
        16'b1111100000011000 : reciprocal = 1111111111111111;
        16'b1111100000010111 : reciprocal = 1111111111111111;
        16'b1111100000010110 : reciprocal = 1111111111111111;
        16'b1111100000010101 : reciprocal = 1111111111111111;
        16'b1111100000010100 : reciprocal = 1111111111111111;
        16'b1111100000010011 : reciprocal = 1111111111111111;
        16'b1111100000010010 : reciprocal = 1111111111111111;
        16'b1111100000010001 : reciprocal = 1111111111111111;
        16'b1111100000010000 : reciprocal = 1111111111111111;
        16'b1111100000001111 : reciprocal = 1111111111111111;
        16'b1111100000001110 : reciprocal = 1111111111111111;
        16'b1111100000001101 : reciprocal = 1111111111111111;
        16'b1111100000001100 : reciprocal = 1111111111111111;
        16'b1111100000001011 : reciprocal = 1111111111111111;
        16'b1111100000001010 : reciprocal = 1111111111111111;
        16'b1111100000001001 : reciprocal = 1111111111111111;
        16'b1111100000001000 : reciprocal = 1111111111111111;
        16'b1111100000000111 : reciprocal = 1111111111111111;
        16'b1111100000000110 : reciprocal = 1111111111111111;
        16'b1111100000000101 : reciprocal = 1111111111111111;
        16'b1111100000000100 : reciprocal = 1111111111111111;
        16'b1111100000000011 : reciprocal = 1111111111111111;
        16'b1111100000000010 : reciprocal = 1111111111111111;
        16'b1111100000000001 : reciprocal = 1111111111111111;


        endcase
    end
    



    //////////////////////// For testbenching ////////////////////////
    // synthesis translate_off

    // synthesis translate_on

endmodule
