// Author: Abdelrahman Elabd
// Lab: ACME Labs, U. Washington ECE
// Date: 04/17/2025
// Module purpose: This module takes an 8bit integer value, 'number_in', and returns a 24-bit fractional value for its reciprocal value, 'reciprocal'. 

module udivision_LUT_8bit_int_to_24bit_frac #(
)(
    input logic [8-1:0] number_in,
    output logic [24-1:0] reciprocal

);

    logic [2**8-1:0] reciprocal_LUT [24-1:0];

    always_comb begin
        case (number_in)
        8'b00000000 : reciprocal = 24'b111111111111111111111111;
        8'b00000001 : reciprocal = 24'b100000000000000000000000;
        8'b00000010 : reciprocal = 24'b010101010101010101010101;
        8'b00000011 : reciprocal = 24'b010000000000000000000000;
        8'b00000100 : reciprocal = 24'b001100110011001100110011;
        8'b00000101 : reciprocal = 24'b001010101010101010101010;
        8'b00000110 : reciprocal = 24'b001001001001001001001001;
        8'b00000111 : reciprocal = 24'b001000000000000000000000;
        8'b00001000 : reciprocal = 24'b000111000111000111000111;
        8'b00001001 : reciprocal = 24'b000110011001100110011001;
        8'b00001010 : reciprocal = 24'b000101110100010111010001;
        8'b00001011 : reciprocal = 24'b000101010101010101010101;
        8'b00001100 : reciprocal = 24'b000100111011000100111011;
        8'b00001101 : reciprocal = 24'b000100100100100100100100;
        8'b00001110 : reciprocal = 24'b000100010001000100010001;
        8'b00001111 : reciprocal = 24'b000100000000000000000000;
        8'b00010000 : reciprocal = 24'b000011110000111100001111;
        8'b00010001 : reciprocal = 24'b000011100011100011100011;
        8'b00010010 : reciprocal = 24'b000011010111100101000011;
        8'b00010011 : reciprocal = 24'b000011001100110011001100;
        8'b00010100 : reciprocal = 24'b000011000011000011000011;
        8'b00010101 : reciprocal = 24'b000010111010001011101000;
        8'b00010110 : reciprocal = 24'b000010110010000101100100;
        8'b00010111 : reciprocal = 24'b000010101010101010101010;
        8'b00011000 : reciprocal = 24'b000010100011110101110000;
        8'b00011001 : reciprocal = 24'b000010011101100010011101;
        8'b00011010 : reciprocal = 24'b000010010111101101000010;
        8'b00011011 : reciprocal = 24'b000010010010010010010010;
        8'b00011100 : reciprocal = 24'b000010001101001111011100;
        8'b00011101 : reciprocal = 24'b000010001000100010001000;
        8'b00011110 : reciprocal = 24'b000010000100001000010000;
        8'b00011111 : reciprocal = 24'b000010000000000000000000;
        8'b00100000 : reciprocal = 24'b000001111100000111110000;
        8'b00100001 : reciprocal = 24'b000001111000011110000111;
        8'b00100010 : reciprocal = 24'b000001110101000001110101;
        8'b00100011 : reciprocal = 24'b000001110001110001110001;
        8'b00100100 : reciprocal = 24'b000001101110101100111110;
        8'b00100101 : reciprocal = 24'b000001101011110010100001;
        8'b00100110 : reciprocal = 24'b000001101001000001101001;
        8'b00100111 : reciprocal = 24'b000001100110011001100110;
        8'b00101000 : reciprocal = 24'b000001100011111001110000;
        8'b00101001 : reciprocal = 24'b000001100001100001100001;
        8'b00101010 : reciprocal = 24'b000001011111010000010111;
        8'b00101011 : reciprocal = 24'b000001011101000101110100;
        8'b00101100 : reciprocal = 24'b000001011011000001011011;
        8'b00101101 : reciprocal = 24'b000001011001000010110010;
        8'b00101110 : reciprocal = 24'b000001010111001001100010;
        8'b00101111 : reciprocal = 24'b000001010101010101010101;
        8'b00110000 : reciprocal = 24'b000001010011100101111000;
        8'b00110001 : reciprocal = 24'b000001010001111010111000;
        8'b00110010 : reciprocal = 24'b000001010000010100000101;
        8'b00110011 : reciprocal = 24'b000001001110110001001110;
        8'b00110100 : reciprocal = 24'b000001001101010010000111;
        8'b00110101 : reciprocal = 24'b000001001011110110100001;
        8'b00110110 : reciprocal = 24'b000001001010011110010000;
        8'b00110111 : reciprocal = 24'b000001001001001001001001;
        8'b00111000 : reciprocal = 24'b000001000111110111000001;
        8'b00111001 : reciprocal = 24'b000001000110100111101110;
        8'b00111010 : reciprocal = 24'b000001000101011011000111;
        8'b00111011 : reciprocal = 24'b000001000100010001000100;
        8'b00111100 : reciprocal = 24'b000001000011001001011100;
        8'b00111101 : reciprocal = 24'b000001000010000100001000;
        8'b00111110 : reciprocal = 24'b000001000001000001000001;
        8'b00111111 : reciprocal = 24'b000001000000000000000000;
        8'b01000000 : reciprocal = 24'b000000111111000000111111;
        8'b01000001 : reciprocal = 24'b000000111110000011111000;
        8'b01000010 : reciprocal = 24'b000000111101001000100110;
        8'b01000011 : reciprocal = 24'b000000111100001111000011;
        8'b01000100 : reciprocal = 24'b000000111011010111001100;
        8'b01000101 : reciprocal = 24'b000000111010100000111010;
        8'b01000110 : reciprocal = 24'b000000111001101100001010;
        8'b01000111 : reciprocal = 24'b000000111000111000111000;
        8'b01001000 : reciprocal = 24'b000000111000000111000000;
        8'b01001001 : reciprocal = 24'b000000110111010110011111;
        8'b01001010 : reciprocal = 24'b000000110110100111010000;
        8'b01001011 : reciprocal = 24'b000000110101111001010000;
        8'b01001100 : reciprocal = 24'b000000110101001100011101;
        8'b01001101 : reciprocal = 24'b000000110100100000110100;
        8'b01001110 : reciprocal = 24'b000000110011110110010001;
        8'b01001111 : reciprocal = 24'b000000110011001100110011;
        8'b01010000 : reciprocal = 24'b000000110010100100010110;
        8'b01010001 : reciprocal = 24'b000000110001111100111000;
        8'b01010010 : reciprocal = 24'b000000110001010110010111;
        8'b01010011 : reciprocal = 24'b000000110000110000110000;
        8'b01010100 : reciprocal = 24'b000000110000001100000011;
        8'b01010101 : reciprocal = 24'b000000101111101000001011;
        8'b01010110 : reciprocal = 24'b000000101111000101001001;
        8'b01010111 : reciprocal = 24'b000000101110100010111010;
        8'b01011000 : reciprocal = 24'b000000101110000001011100;
        8'b01011001 : reciprocal = 24'b000000101101100000101101;
        8'b01011010 : reciprocal = 24'b000000101101000000101101;
        8'b01011011 : reciprocal = 24'b000000101100100001011001;
        8'b01011100 : reciprocal = 24'b000000101100000010110000;
        8'b01011101 : reciprocal = 24'b000000101011100100110001;
        8'b01011110 : reciprocal = 24'b000000101011000111011010;
        8'b01011111 : reciprocal = 24'b000000101010101010101010;
        8'b01100000 : reciprocal = 24'b000000101010001110100000;
        8'b01100001 : reciprocal = 24'b000000101001110010111100;
        8'b01100010 : reciprocal = 24'b000000101001010111111010;
        8'b01100011 : reciprocal = 24'b000000101000111101011100;
        8'b01100100 : reciprocal = 24'b000000101000100011011111;
        8'b01100101 : reciprocal = 24'b000000101000001010000010;
        8'b01100110 : reciprocal = 24'b000000100111110001000101;
        8'b01100111 : reciprocal = 24'b000000100111011000100111;
        8'b01101000 : reciprocal = 24'b000000100111000000100111;
        8'b01101001 : reciprocal = 24'b000000100110101001000011;
        8'b01101010 : reciprocal = 24'b000000100110010001111100;
        8'b01101011 : reciprocal = 24'b000000100101111011010000;
        8'b01101100 : reciprocal = 24'b000000100101100100111111;
        8'b01101101 : reciprocal = 24'b000000100101001111001000;
        8'b01101110 : reciprocal = 24'b000000100100111001101010;
        8'b01101111 : reciprocal = 24'b000000100100100100100100;
        8'b01110000 : reciprocal = 24'b000000100100001111110110;
        8'b01110001 : reciprocal = 24'b000000100011111011100000;
        8'b01110010 : reciprocal = 24'b000000100011100111100000;
        8'b01110011 : reciprocal = 24'b000000100011010011110111;
        8'b01110100 : reciprocal = 24'b000000100011000000100011;
        8'b01110101 : reciprocal = 24'b000000100010101101100011;
        8'b01110110 : reciprocal = 24'b000000100010011010111001;
        8'b01110111 : reciprocal = 24'b000000100010001000100010;
        8'b01111000 : reciprocal = 24'b000000100001110110011110;
        8'b01111001 : reciprocal = 24'b000000100001100100101110;
        8'b01111010 : reciprocal = 24'b000000100001010011010000;
        8'b01111011 : reciprocal = 24'b000000100001000010000100;
        8'b01111100 : reciprocal = 24'b000000100000110001001001;
        8'b01111101 : reciprocal = 24'b000000100000100000100000;
        8'b01111110 : reciprocal = 24'b000000100000010000001000;
        8'b01111111 : reciprocal = 24'b000000100000000000000000;
        8'b10000000 : reciprocal = 24'b000000011111110000000111;
        8'b10000001 : reciprocal = 24'b000000011111100000011111;
        8'b10000010 : reciprocal = 24'b000000011111010001000110;
        8'b10000011 : reciprocal = 24'b000000011111000001111100;
        8'b10000100 : reciprocal = 24'b000000011110110011000000;
        8'b10000101 : reciprocal = 24'b000000011110100100010011;
        8'b10000110 : reciprocal = 24'b000000011110010101110011;
        8'b10000111 : reciprocal = 24'b000000011110000111100001;
        8'b10001000 : reciprocal = 24'b000000011101111001011101;
        8'b10001001 : reciprocal = 24'b000000011101101011100110;
        8'b10001010 : reciprocal = 24'b000000011101011101111011;
        8'b10001011 : reciprocal = 24'b000000011101010000011101;
        8'b10001100 : reciprocal = 24'b000000011101000011001011;
        8'b10001101 : reciprocal = 24'b000000011100110110000101;
        8'b10001110 : reciprocal = 24'b000000011100101001001011;
        8'b10001111 : reciprocal = 24'b000000011100011100011100;
        8'b10010000 : reciprocal = 24'b000000011100001111111000;
        8'b10010001 : reciprocal = 24'b000000011100000011100000;
        8'b10010010 : reciprocal = 24'b000000011011110111010010;
        8'b10010011 : reciprocal = 24'b000000011011101011001111;
        8'b10010100 : reciprocal = 24'b000000011011011111010110;
        8'b10010101 : reciprocal = 24'b000000011011010011101000;
        8'b10010110 : reciprocal = 24'b000000011011001000000011;
        8'b10010111 : reciprocal = 24'b000000011010111100101000;
        8'b10011000 : reciprocal = 24'b000000011010110001010111;
        8'b10011001 : reciprocal = 24'b000000011010100110001110;
        8'b10011010 : reciprocal = 24'b000000011010011011010000;
        8'b10011011 : reciprocal = 24'b000000011010010000011010;
        8'b10011100 : reciprocal = 24'b000000011010000101101101;
        8'b10011101 : reciprocal = 24'b000000011001111011001000;
        8'b10011110 : reciprocal = 24'b000000011001110000101101;
        8'b10011111 : reciprocal = 24'b000000011001100110011001;
        8'b10100000 : reciprocal = 24'b000000011001011100001110;
        8'b10100001 : reciprocal = 24'b000000011001010010001011;
        8'b10100010 : reciprocal = 24'b000000011001001000001111;
        8'b10100011 : reciprocal = 24'b000000011000111110011100;
        8'b10100100 : reciprocal = 24'b000000011000110100110000;
        8'b10100101 : reciprocal = 24'b000000011000101011001011;
        8'b10100110 : reciprocal = 24'b000000011000100001101110;
        8'b10100111 : reciprocal = 24'b000000011000011000011000;
        8'b10101000 : reciprocal = 24'b000000011000001111001001;
        8'b10101001 : reciprocal = 24'b000000011000000110000001;
        8'b10101010 : reciprocal = 24'b000000010111111101000000;
        8'b10101011 : reciprocal = 24'b000000010111110100000101;
        8'b10101100 : reciprocal = 24'b000000010111101011010010;
        8'b10101101 : reciprocal = 24'b000000010111100010100100;
        8'b10101110 : reciprocal = 24'b000000010111011001111101;
        8'b10101111 : reciprocal = 24'b000000010111010001011101;
        8'b10110000 : reciprocal = 24'b000000010111001001000010;
        8'b10110001 : reciprocal = 24'b000000010111000000101110;
        8'b10110010 : reciprocal = 24'b000000010110111000011111;
        8'b10110011 : reciprocal = 24'b000000010110110000010110;
        8'b10110100 : reciprocal = 24'b000000010110101000010011;
        8'b10110101 : reciprocal = 24'b000000010110100000010110;
        8'b10110110 : reciprocal = 24'b000000010110011000011110;
        8'b10110111 : reciprocal = 24'b000000010110010000101100;
        8'b10111000 : reciprocal = 24'b000000010110001000111111;
        8'b10111001 : reciprocal = 24'b000000010110000001011000;
        8'b10111010 : reciprocal = 24'b000000010101111001110101;
        8'b10111011 : reciprocal = 24'b000000010101110010011000;
        8'b10111100 : reciprocal = 24'b000000010101101011000000;
        8'b10111101 : reciprocal = 24'b000000010101100011101101;
        8'b10111110 : reciprocal = 24'b000000010101011100011110;
        8'b10111111 : reciprocal = 24'b000000010101010101010101;
        8'b11000000 : reciprocal = 24'b000000010101001110010000;
        8'b11000001 : reciprocal = 24'b000000010101000111010000;
        8'b11000010 : reciprocal = 24'b000000010101000000010101;
        8'b11000011 : reciprocal = 24'b000000010100111001011110;
        8'b11000100 : reciprocal = 24'b000000010100110010101011;
        8'b11000101 : reciprocal = 24'b000000010100101011111101;
        8'b11000110 : reciprocal = 24'b000000010100100101010011;
        8'b11000111 : reciprocal = 24'b000000010100011110101110;
        8'b11001000 : reciprocal = 24'b000000010100011000001100;
        8'b11001001 : reciprocal = 24'b000000010100010001101111;
        8'b11001010 : reciprocal = 24'b000000010100001011010110;
        8'b11001011 : reciprocal = 24'b000000010100000101000001;
        8'b11001100 : reciprocal = 24'b000000010011111110110000;
        8'b11001101 : reciprocal = 24'b000000010011111000100010;
        8'b11001110 : reciprocal = 24'b000000010011110010011001;
        8'b11001111 : reciprocal = 24'b000000010011101100010011;
        8'b11010000 : reciprocal = 24'b000000010011100110010001;
        8'b11010001 : reciprocal = 24'b000000010011100000010011;
        8'b11010010 : reciprocal = 24'b000000010011011010011000;
        8'b11010011 : reciprocal = 24'b000000010011010100100001;
        8'b11010100 : reciprocal = 24'b000000010011001110101110;
        8'b11010101 : reciprocal = 24'b000000010011001000111110;
        8'b11010110 : reciprocal = 24'b000000010011000011010001;
        8'b11010111 : reciprocal = 24'b000000010010111101101000;
        8'b11011000 : reciprocal = 24'b000000010010111000000010;
        8'b11011001 : reciprocal = 24'b000000010010110010011111;
        8'b11011010 : reciprocal = 24'b000000010010101101000000;
        8'b11011011 : reciprocal = 24'b000000010010100111100100;
        8'b11011100 : reciprocal = 24'b000000010010100010001011;
        8'b11011101 : reciprocal = 24'b000000010010011100110101;
        8'b11011110 : reciprocal = 24'b000000010010010111100010;
        8'b11011111 : reciprocal = 24'b000000010010010010010010;
        8'b11100000 : reciprocal = 24'b000000010010001101000101;
        8'b11100001 : reciprocal = 24'b000000010010000111111011;
        8'b11100010 : reciprocal = 24'b000000010010000010110100;
        8'b11100011 : reciprocal = 24'b000000010001111101110000;
        8'b11100100 : reciprocal = 24'b000000010001111000101110;
        8'b11100101 : reciprocal = 24'b000000010001110011110000;
        8'b11100110 : reciprocal = 24'b000000010001101110110100;
        8'b11100111 : reciprocal = 24'b000000010001101001111011;
        8'b11101000 : reciprocal = 24'b000000010001100101000101;
        8'b11101001 : reciprocal = 24'b000000010001100000010001;
        8'b11101010 : reciprocal = 24'b000000010001011011100000;
        8'b11101011 : reciprocal = 24'b000000010001010110110001;
        8'b11101100 : reciprocal = 24'b000000010001010010000101;
        8'b11101101 : reciprocal = 24'b000000010001001101011100;
        8'b11101110 : reciprocal = 24'b000000010001001000110101;
        8'b11101111 : reciprocal = 24'b000000010001000100010001;
        8'b11110000 : reciprocal = 24'b000000010000111111101111;
        8'b11110001 : reciprocal = 24'b000000010000111011001111;
        8'b11110010 : reciprocal = 24'b000000010000110110110010;
        8'b11110011 : reciprocal = 24'b000000010000110010010111;
        8'b11110100 : reciprocal = 24'b000000010000101101111110;
        8'b11110101 : reciprocal = 24'b000000010000101001101000;
        8'b11110110 : reciprocal = 24'b000000010000100101010011;
        8'b11110111 : reciprocal = 24'b000000010000100001000010;
        8'b11111000 : reciprocal = 24'b000000010000011100110010;
        8'b11111001 : reciprocal = 24'b000000010000011000100100;
        8'b11111010 : reciprocal = 24'b000000010000010100011001;
        8'b11111011 : reciprocal = 24'b000000010000010000010000;
        8'b11111100 : reciprocal = 24'b000000010000001100001001;
        8'b11111101 : reciprocal = 24'b000000010000001000000100;
        8'b11111110 : reciprocal = 24'b000000010000000100000001;
        8'b11111111 : reciprocal = 24'b000000010000000000000000;


        endcase
    end
    



    //////////////////////// For testbenching ////////////////////////
    // synthesis translate_off

    // synthesis translate_on

endmodule
