module norm_reader #(
    parameter PIXEL_BIT_WIDTH   = 10,
    parameter OUT_ROWS          = 10,
    parameter OUT_COLS          = 10
)(
    input  logic                     clk,
    input  logic                     srst,
    input  logic                     s_axis_resetn,

    // ap control signals
    input logic seq_ap_idle,
    input logic cf_ap_done,

    input logic ap_start, 
    output logic ap_done,
    output logic ap_ready, 
    // output logic ap_idle, // TODO

    // AXI Stream Slave Interface
    input  logic                     s_axis_tvalid,
    output logic                     s_axis_tready,
    input  logic [PIXEL_BIT_WIDTH-1:0] s_axis_tdata,

    // Normalization value
    input logic [PIXEL_BIT_WIDTH-1:0] norm_denominator,

    // AXI Stream Master Interface
    output logic                   m_axis_tvalid,
    input  logic                   m_axis_tready,
    output logic [PIXEL_BIT_WIDTH-1:0] m_axis_tdata

);

    logic intmd_axis_tvalid;
    logic intmd_axis_tready;
    logic [PIXEL_BIT_WIDTH-1:0] intmd_axis_tdata;

    axis_fifo nr_axis_fifo (.s_aclk(clk),
                            .s_aresetn(~reset),
                            .s_axis_tvalid(intmd_axis_tvalid),
                            .s_axis_tready(intmd_axis_tready),
                            .s_axis_tdata(intmd_axis_tdata),
                            .m_axis_tvalid(m_axis_tvalid),
                            .m_axis_tready(m_axis_tready),
                            .m_axis_tdata(m_axis_tdata)
                            );


    // Combine both reset signals into one for simplicity
    logic reset;
    assign reset = srst || (!s_axis_resetn);

    
    //////////////////////// ap_ready ////////////////////////
    logic [$clog2(OUT_ROWS*OUT_COLS)-1:0] cnt_fifo_reads;
    always_ff @(posedge clk) begin
        if (reset || ap_start) cnt_fifo_reads <= 0;
        else if (cnt_fifo_reads == OUT_ROWS*OUT_COLS-1) cnt_fifo_reads <= 0;
        else if (m_axis_tvalid && m_axis_tready) cnt_fifo_reads <= cnt_fifo_reads + 1;
    end

    enum logic {IDLE, NORMALIZING} ps, ns;
    always_ff @(posedge clk) begin
        if (reset) ps <= IDLE;
        else ps <= ns;
    end
    always_comb begin
        case(ps)
            IDLE: begin
                ap_ready = 1'b1;
                if (ap_start && seq_ap_idle) ns = NORMALIZING;
                else ns = IDLE;
            end
            NORMALIZING: begin
                ap_ready = 1'b0;
                if (cnt_fifo_reads == OUT_ROWS*OUT_COLS-1) ns = IDLE;
                else ns = NORMALIZING;
            end
        endcase
    end

    //////////////////////// ready_to_norm: only true if the upstream crop-filter is done with its task ////////////////////////
    logic ready_to_norm;
    always_ff @(posedge clk) begin
        if (reset || ap_start) begin
            ready_to_norm <= 1'b0;
        end
        else if (cf_ap_done) begin
            ready_to_norm <= 1'b1;
        end
    end 


    //////////////////////// Normalization logic ////////////////////////

    // reciprocal of max value to get normalization coefficient
    logic [PIXEL_BIT_WIDTH-1:0] norm_coef;
    udivision_LUT_8bit_int_to_8bit_frac norm_coef_getter (.number_in(norm_denominator), .reciprocal(norm_coef));

    // multiplication: 
    umult_int_frac #(.WIDTH(PIXEL_BIT_WIDTH)) normed_pixel_getter (.pixel(s_axis_tdata), .norm_factor(norm_coef), .out(intmd_axis_tdata));
    // assign intmd_axis_tdata = s_axis_tdata; 

    // assign s_axis_tready = ready_to_norm && m_axis_tready;
    assign s_axis_tready = intmd_axis_tready && ready_to_norm; // pass-through for now
    assign intmd_axis_tvalid = s_axis_tvalid && ready_to_norm;
    
    
    //////////////////////// For testbenching ////////////////////////
    // synthesis translate_off

    // synthesis translate_on

endmodule
